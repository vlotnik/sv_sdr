    DVBS2_BPSK : super.plane = {
           0.707    ,  0.707            // 0
        , -0.707    , -0.707            // 1
    };