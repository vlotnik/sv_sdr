    QAM2048 : super.plane = {
           2.747    ,  2.924            // 0
        ,  2.569    ,  2.924            // 1
        ,  2.747    ,  3.101            // 2
        ,  2.569    ,  3.101            // 3
        ,  2.215    ,  2.924            // 4
        ,  2.392    ,  2.924            // 5
        ,  2.215    ,  3.101            // 6
        ,  2.392    ,  3.101            // 7
        ,  2.747    ,  3.455            // 8
        ,  2.569    ,  3.455            // 9
        ,  2.747    ,  3.278            // 10
        ,  2.569    ,  3.278            // 11
        ,  2.215    ,  3.455            // 12
        ,  2.392    ,  3.455            // 13
        ,  2.215    ,  3.278            // 14
        ,  2.392    ,  3.278            // 15
        ,  1.506    ,  2.924            // 16
        ,  1.683    ,  2.924            // 17
        ,  1.506    ,  3.101            // 18
        ,  1.683    ,  3.101            // 19
        ,  2.038    ,  2.924            // 20
        ,  1.861    ,  2.924            // 21
        ,  2.038    ,  3.101            // 22
        ,  1.861    ,  3.101            // 23
        ,  1.506    ,  3.455            // 24
        ,  1.683    ,  3.455            // 25
        ,  1.506    ,  3.278            // 26
        ,  1.683    ,  3.278            // 27
        ,  2.038    ,  3.455            // 28
        ,  1.861    ,  3.455            // 29
        ,  2.038    ,  3.278            // 30
        ,  1.861    ,  3.278            // 31
        ,  2.747    ,  4.164            // 32
        ,  2.569    ,  4.164            // 33
        ,  2.747    ,  3.987            // 34
        ,  2.569    ,  3.987            // 35
        ,  2.215    ,  4.164            // 36
        ,  2.392    ,  4.164            // 37
        ,  2.215    ,  3.987            // 38
        ,  2.392    ,  3.987            // 39
        ,  2.747    ,  3.633            // 40
        ,  2.569    ,  3.633            // 41
        ,  2.747    ,   3.81            // 42
        ,  2.569    ,   3.81            // 43
        ,  2.215    ,  3.633            // 44
        ,  2.392    ,  3.633            // 45
        ,  2.215    ,   3.81            // 46
        ,  2.392    ,   3.81            // 47
        ,  1.506    ,  4.164            // 48
        ,  1.683    ,  4.164            // 49
        ,  1.506    ,  3.987            // 50
        ,  1.683    ,  3.987            // 51
        ,  2.038    ,  4.164            // 52
        ,  1.861    ,  4.164            // 53
        ,  2.038    ,  3.987            // 54
        ,  1.861    ,  3.987            // 55
        ,  1.506    ,  3.633            // 56
        ,  1.683    ,  3.633            // 57
        ,  1.506    ,   3.81            // 58
        ,  1.683    ,   3.81            // 59
        ,  2.038    ,  3.633            // 60
        ,  1.861    ,  3.633            // 61
        ,  2.038    ,   3.81            // 62
        ,  1.861    ,   3.81            // 63
        ,  2.924    ,  2.747            // 64
        ,  3.101    ,  2.747            // 65
        ,  2.924    ,  2.569            // 66
        ,  3.101    ,  2.569            // 67
        ,  3.455    ,  2.747            // 68
        ,  3.278    ,  2.747            // 69
        ,  3.455    ,  2.569            // 70
        ,  3.278    ,  2.569            // 71
        ,  2.924    ,  2.215            // 72
        ,  3.101    ,  2.215            // 73
        ,  2.924    ,  2.392            // 74
        ,  3.101    ,  2.392            // 75
        ,  3.455    ,  2.215            // 76
        ,  3.278    ,  2.215            // 77
        ,  3.455    ,  2.392            // 78
        ,  3.278    ,  2.392            // 79
        ,  4.164    ,  2.747            // 80
        ,  3.987    ,  2.747            // 81
        ,  4.164    ,  2.569            // 82
        ,  3.987    ,  2.569            // 83
        ,  3.633    ,  2.747            // 84
        ,   3.81    ,  2.747            // 85
        ,  3.633    ,  2.569            // 86
        ,   3.81    ,  2.569            // 87
        ,  4.164    ,  2.215            // 88
        ,  3.987    ,  2.215            // 89
        ,  4.164    ,  2.392            // 90
        ,  3.987    ,  2.392            // 91
        ,  3.633    ,  2.215            // 92
        ,   3.81    ,  2.215            // 93
        ,  3.633    ,  2.392            // 94
        ,   3.81    ,  2.392            // 95
        ,  2.924    ,  1.506            // 96
        ,  3.101    ,  1.506            // 97
        ,  2.924    ,  1.683            // 98
        ,  3.101    ,  1.683            // 99
        ,  3.455    ,  1.506            // 100
        ,  3.278    ,  1.506            // 101
        ,  3.455    ,  1.683            // 102
        ,  3.278    ,  1.683            // 103
        ,  2.924    ,  2.038            // 104
        ,  3.101    ,  2.038            // 105
        ,  2.924    ,  1.861            // 106
        ,  3.101    ,  1.861            // 107
        ,  3.455    ,  2.038            // 108
        ,  3.278    ,  2.038            // 109
        ,  3.455    ,  1.861            // 110
        ,  3.278    ,  1.861            // 111
        ,  4.164    ,  1.506            // 112
        ,  3.987    ,  1.506            // 113
        ,  4.164    ,  1.683            // 114
        ,  3.987    ,  1.683            // 115
        ,  3.633    ,  1.506            // 116
        ,   3.81    ,  1.506            // 117
        ,  3.633    ,  1.683            // 118
        ,   3.81    ,  1.683            // 119
        ,  4.164    ,  2.038            // 120
        ,  3.987    ,  2.038            // 121
        ,  4.164    ,  1.861            // 122
        ,  3.987    ,  1.861            // 123
        ,  3.633    ,  2.038            // 124
        ,   3.81    ,  2.038            // 125
        ,  3.633    ,  1.861            // 126
        ,   3.81    ,  1.861            // 127
        ,  0.089    ,  2.924            // 128
        ,  0.266    ,  2.924            // 129
        ,  0.089    ,  3.101            // 130
        ,  0.266    ,  3.101            // 131
        ,   0.62    ,  2.924            // 132
        ,  0.443    ,  2.924            // 133
        ,   0.62    ,  3.101            // 134
        ,  0.443    ,  3.101            // 135
        ,  0.089    ,  3.455            // 136
        ,  0.266    ,  3.455            // 137
        ,  0.089    ,  3.278            // 138
        ,  0.266    ,  3.278            // 139
        ,   0.62    ,  3.455            // 140
        ,  0.443    ,  3.455            // 141
        ,   0.62    ,  3.278            // 142
        ,  0.443    ,  3.278            // 143
        ,  1.329    ,  2.924            // 144
        ,  1.152    ,  2.924            // 145
        ,  1.329    ,  3.101            // 146
        ,  1.152    ,  3.101            // 147
        ,  0.797    ,  2.924            // 148
        ,  0.975    ,  2.924            // 149
        ,  0.797    ,  3.101            // 150
        ,  0.975    ,  3.101            // 151
        ,  1.329    ,  3.455            // 152
        ,  1.152    ,  3.455            // 153
        ,  1.329    ,  3.278            // 154
        ,  1.152    ,  3.278            // 155
        ,  0.797    ,  3.455            // 156
        ,  0.975    ,  3.455            // 157
        ,  0.797    ,  3.278            // 158
        ,  0.975    ,  3.278            // 159
        ,  0.089    ,  4.164            // 160
        ,  0.266    ,  4.164            // 161
        ,  0.089    ,  3.987            // 162
        ,  0.266    ,  3.987            // 163
        ,   0.62    ,  4.164            // 164
        ,  0.443    ,  4.164            // 165
        ,   0.62    ,  3.987            // 166
        ,  0.443    ,  3.987            // 167
        ,  0.089    ,  3.633            // 168
        ,  0.266    ,  3.633            // 169
        ,  0.089    ,   3.81            // 170
        ,  0.266    ,   3.81            // 171
        ,   0.62    ,  3.633            // 172
        ,  0.443    ,  3.633            // 173
        ,   0.62    ,   3.81            // 174
        ,  0.443    ,   3.81            // 175
        ,  1.329    ,  4.164            // 176
        ,  1.152    ,  4.164            // 177
        ,  1.329    ,  3.987            // 178
        ,  1.152    ,  3.987            // 179
        ,  0.797    ,  4.164            // 180
        ,  0.975    ,  4.164            // 181
        ,  0.797    ,  3.987            // 182
        ,  0.975    ,  3.987            // 183
        ,  1.329    ,  3.633            // 184
        ,  1.152    ,  3.633            // 185
        ,  1.329    ,   3.81            // 186
        ,  1.152    ,   3.81            // 187
        ,  0.797    ,  3.633            // 188
        ,  0.975    ,  3.633            // 189
        ,  0.797    ,   3.81            // 190
        ,  0.975    ,   3.81            // 191
        ,  2.924    ,  0.089            // 192
        ,  3.101    ,  0.089            // 193
        ,  2.924    ,  0.266            // 194
        ,  3.101    ,  0.266            // 195
        ,  3.455    ,  0.089            // 196
        ,  3.278    ,  0.089            // 197
        ,  3.455    ,  0.266            // 198
        ,  3.278    ,  0.266            // 199
        ,  2.924    ,   0.62            // 200
        ,  3.101    ,   0.62            // 201
        ,  2.924    ,  0.443            // 202
        ,  3.101    ,  0.443            // 203
        ,  3.455    ,   0.62            // 204
        ,  3.278    ,   0.62            // 205
        ,  3.455    ,  0.443            // 206
        ,  3.278    ,  0.443            // 207
        ,  4.164    ,  0.089            // 208
        ,  3.987    ,  0.089            // 209
        ,  4.164    ,  0.266            // 210
        ,  3.987    ,  0.266            // 211
        ,  3.633    ,  0.089            // 212
        ,   3.81    ,  0.089            // 213
        ,  3.633    ,  0.266            // 214
        ,   3.81    ,  0.266            // 215
        ,  4.164    ,   0.62            // 216
        ,  3.987    ,   0.62            // 217
        ,  4.164    ,  0.443            // 218
        ,  3.987    ,  0.443            // 219
        ,  3.633    ,   0.62            // 220
        ,   3.81    ,   0.62            // 221
        ,  3.633    ,  0.443            // 222
        ,   3.81    ,  0.443            // 223
        ,  2.924    ,  1.329            // 224
        ,  3.101    ,  1.329            // 225
        ,  2.924    ,  1.152            // 226
        ,  3.101    ,  1.152            // 227
        ,  3.455    ,  1.329            // 228
        ,  3.278    ,  1.329            // 229
        ,  3.455    ,  1.152            // 230
        ,  3.278    ,  1.152            // 231
        ,  2.924    ,  0.797            // 232
        ,  3.101    ,  0.797            // 233
        ,  2.924    ,  0.975            // 234
        ,  3.101    ,  0.975            // 235
        ,  3.455    ,  0.797            // 236
        ,  3.278    ,  0.797            // 237
        ,  3.455    ,  0.975            // 238
        ,  3.278    ,  0.975            // 239
        ,  4.164    ,  1.329            // 240
        ,  3.987    ,  1.329            // 241
        ,  4.164    ,  1.152            // 242
        ,  3.987    ,  1.152            // 243
        ,  3.633    ,  1.329            // 244
        ,   3.81    ,  1.329            // 245
        ,  3.633    ,  1.152            // 246
        ,   3.81    ,  1.152            // 247
        ,  4.164    ,  0.797            // 248
        ,  3.987    ,  0.797            // 249
        ,  4.164    ,  0.975            // 250
        ,  3.987    ,  0.975            // 251
        ,  3.633    ,  0.797            // 252
        ,   3.81    ,  0.797            // 253
        ,  3.633    ,  0.975            // 254
        ,   3.81    ,  0.975            // 255
        ,  0.089    ,  2.747            // 256
        ,  0.266    ,  2.747            // 257
        ,  0.089    ,  2.569            // 258
        ,  0.266    ,  2.569            // 259
        ,   0.62    ,  2.747            // 260
        ,  0.443    ,  2.747            // 261
        ,   0.62    ,  2.569            // 262
        ,  0.443    ,  2.569            // 263
        ,  0.089    ,  2.215            // 264
        ,  0.266    ,  2.215            // 265
        ,  0.089    ,  2.392            // 266
        ,  0.266    ,  2.392            // 267
        ,   0.62    ,  2.215            // 268
        ,  0.443    ,  2.215            // 269
        ,   0.62    ,  2.392            // 270
        ,  0.443    ,  2.392            // 271
        ,  1.329    ,  2.747            // 272
        ,  1.152    ,  2.747            // 273
        ,  1.329    ,  2.569            // 274
        ,  1.152    ,  2.569            // 275
        ,  0.797    ,  2.747            // 276
        ,  0.975    ,  2.747            // 277
        ,  0.797    ,  2.569            // 278
        ,  0.975    ,  2.569            // 279
        ,  1.329    ,  2.215            // 280
        ,  1.152    ,  2.215            // 281
        ,  1.329    ,  2.392            // 282
        ,  1.152    ,  2.392            // 283
        ,  0.797    ,  2.215            // 284
        ,  0.975    ,  2.215            // 285
        ,  0.797    ,  2.392            // 286
        ,  0.975    ,  2.392            // 287
        ,  0.089    ,  1.506            // 288
        ,  0.266    ,  1.506            // 289
        ,  0.089    ,  1.683            // 290
        ,  0.266    ,  1.683            // 291
        ,   0.62    ,  1.506            // 292
        ,  0.443    ,  1.506            // 293
        ,   0.62    ,  1.683            // 294
        ,  0.443    ,  1.683            // 295
        ,  0.089    ,  2.038            // 296
        ,  0.266    ,  2.038            // 297
        ,  0.089    ,  1.861            // 298
        ,  0.266    ,  1.861            // 299
        ,   0.62    ,  2.038            // 300
        ,  0.443    ,  2.038            // 301
        ,   0.62    ,  1.861            // 302
        ,  0.443    ,  1.861            // 303
        ,  1.329    ,  1.506            // 304
        ,  1.152    ,  1.506            // 305
        ,  1.329    ,  1.683            // 306
        ,  1.152    ,  1.683            // 307
        ,  0.797    ,  1.506            // 308
        ,  0.975    ,  1.506            // 309
        ,  0.797    ,  1.683            // 310
        ,  0.975    ,  1.683            // 311
        ,  1.329    ,  2.038            // 312
        ,  1.152    ,  2.038            // 313
        ,  1.329    ,  1.861            // 314
        ,  1.152    ,  1.861            // 315
        ,  0.797    ,  2.038            // 316
        ,  0.975    ,  2.038            // 317
        ,  0.797    ,  1.861            // 318
        ,  0.975    ,  1.861            // 319
        ,  2.747    ,  2.747            // 320
        ,  2.569    ,  2.747            // 321
        ,  2.747    ,  2.569            // 322
        ,  2.569    ,  2.569            // 323
        ,  2.215    ,  2.747            // 324
        ,  2.392    ,  2.747            // 325
        ,  2.215    ,  2.569            // 326
        ,  2.392    ,  2.569            // 327
        ,  2.747    ,  2.215            // 328
        ,  2.569    ,  2.215            // 329
        ,  2.747    ,  2.392            // 330
        ,  2.569    ,  2.392            // 331
        ,  2.215    ,  2.215            // 332
        ,  2.392    ,  2.215            // 333
        ,  2.215    ,  2.392            // 334
        ,  2.392    ,  2.392            // 335
        ,  1.506    ,  2.747            // 336
        ,  1.683    ,  2.747            // 337
        ,  1.506    ,  2.569            // 338
        ,  1.683    ,  2.569            // 339
        ,  2.038    ,  2.747            // 340
        ,  1.861    ,  2.747            // 341
        ,  2.038    ,  2.569            // 342
        ,  1.861    ,  2.569            // 343
        ,  1.506    ,  2.215            // 344
        ,  1.683    ,  2.215            // 345
        ,  1.506    ,  2.392            // 346
        ,  1.683    ,  2.392            // 347
        ,  2.038    ,  2.215            // 348
        ,  1.861    ,  2.215            // 349
        ,  2.038    ,  2.392            // 350
        ,  1.861    ,  2.392            // 351
        ,  2.747    ,  1.506            // 352
        ,  2.569    ,  1.506            // 353
        ,  2.747    ,  1.683            // 354
        ,  2.569    ,  1.683            // 355
        ,  2.215    ,  1.506            // 356
        ,  2.392    ,  1.506            // 357
        ,  2.215    ,  1.683            // 358
        ,  2.392    ,  1.683            // 359
        ,  2.747    ,  2.038            // 360
        ,  2.569    ,  2.038            // 361
        ,  2.747    ,  1.861            // 362
        ,  2.569    ,  1.861            // 363
        ,  2.215    ,  2.038            // 364
        ,  2.392    ,  2.038            // 365
        ,  2.215    ,  1.861            // 366
        ,  2.392    ,  1.861            // 367
        ,  1.506    ,  1.506            // 368
        ,  1.683    ,  1.506            // 369
        ,  1.506    ,  1.683            // 370
        ,  1.683    ,  1.683            // 371
        ,  2.038    ,  1.506            // 372
        ,  1.861    ,  1.506            // 373
        ,  2.038    ,  1.683            // 374
        ,  1.861    ,  1.683            // 375
        ,  1.506    ,  2.038            // 376
        ,  1.683    ,  2.038            // 377
        ,  1.506    ,  1.861            // 378
        ,  1.683    ,  1.861            // 379
        ,  2.038    ,  2.038            // 380
        ,  1.861    ,  2.038            // 381
        ,  2.038    ,  1.861            // 382
        ,  1.861    ,  1.861            // 383
        ,  0.089    ,  0.089            // 384
        ,  0.266    ,  0.089            // 385
        ,  0.089    ,  0.266            // 386
        ,  0.266    ,  0.266            // 387
        ,   0.62    ,  0.089            // 388
        ,  0.443    ,  0.089            // 389
        ,   0.62    ,  0.266            // 390
        ,  0.443    ,  0.266            // 391
        ,  0.089    ,   0.62            // 392
        ,  0.266    ,   0.62            // 393
        ,  0.089    ,  0.443            // 394
        ,  0.266    ,  0.443            // 395
        ,   0.62    ,   0.62            // 396
        ,  0.443    ,   0.62            // 397
        ,   0.62    ,  0.443            // 398
        ,  0.443    ,  0.443            // 399
        ,  1.329    ,  0.089            // 400
        ,  1.152    ,  0.089            // 401
        ,  1.329    ,  0.266            // 402
        ,  1.152    ,  0.266            // 403
        ,  0.797    ,  0.089            // 404
        ,  0.975    ,  0.089            // 405
        ,  0.797    ,  0.266            // 406
        ,  0.975    ,  0.266            // 407
        ,  1.329    ,   0.62            // 408
        ,  1.152    ,   0.62            // 409
        ,  1.329    ,  0.443            // 410
        ,  1.152    ,  0.443            // 411
        ,  0.797    ,   0.62            // 412
        ,  0.975    ,   0.62            // 413
        ,  0.797    ,  0.443            // 414
        ,  0.975    ,  0.443            // 415
        ,  0.089    ,  1.329            // 416
        ,  0.266    ,  1.329            // 417
        ,  0.089    ,  1.152            // 418
        ,  0.266    ,  1.152            // 419
        ,   0.62    ,  1.329            // 420
        ,  0.443    ,  1.329            // 421
        ,   0.62    ,  1.152            // 422
        ,  0.443    ,  1.152            // 423
        ,  0.089    ,  0.797            // 424
        ,  0.266    ,  0.797            // 425
        ,  0.089    ,  0.975            // 426
        ,  0.266    ,  0.975            // 427
        ,   0.62    ,  0.797            // 428
        ,  0.443    ,  0.797            // 429
        ,   0.62    ,  0.975            // 430
        ,  0.443    ,  0.975            // 431
        ,  1.329    ,  1.329            // 432
        ,  1.152    ,  1.329            // 433
        ,  1.329    ,  1.152            // 434
        ,  1.152    ,  1.152            // 435
        ,  0.797    ,  1.329            // 436
        ,  0.975    ,  1.329            // 437
        ,  0.797    ,  1.152            // 438
        ,  0.975    ,  1.152            // 439
        ,  1.329    ,  0.797            // 440
        ,  1.152    ,  0.797            // 441
        ,  1.329    ,  0.975            // 442
        ,  1.152    ,  0.975            // 443
        ,  0.797    ,  0.797            // 444
        ,  0.975    ,  0.797            // 445
        ,  0.797    ,  0.975            // 446
        ,  0.975    ,  0.975            // 447
        ,  2.747    ,  0.089            // 448
        ,  2.569    ,  0.089            // 449
        ,  2.747    ,  0.266            // 450
        ,  2.569    ,  0.266            // 451
        ,  2.215    ,  0.089            // 452
        ,  2.392    ,  0.089            // 453
        ,  2.215    ,  0.266            // 454
        ,  2.392    ,  0.266            // 455
        ,  2.747    ,   0.62            // 456
        ,  2.569    ,   0.62            // 457
        ,  2.747    ,  0.443            // 458
        ,  2.569    ,  0.443            // 459
        ,  2.215    ,   0.62            // 460
        ,  2.392    ,   0.62            // 461
        ,  2.215    ,  0.443            // 462
        ,  2.392    ,  0.443            // 463
        ,  1.506    ,  0.089            // 464
        ,  1.683    ,  0.089            // 465
        ,  1.506    ,  0.266            // 466
        ,  1.683    ,  0.266            // 467
        ,  2.038    ,  0.089            // 468
        ,  1.861    ,  0.089            // 469
        ,  2.038    ,  0.266            // 470
        ,  1.861    ,  0.266            // 471
        ,  1.506    ,   0.62            // 472
        ,  1.683    ,   0.62            // 473
        ,  1.506    ,  0.443            // 474
        ,  1.683    ,  0.443            // 475
        ,  2.038    ,   0.62            // 476
        ,  1.861    ,   0.62            // 477
        ,  2.038    ,  0.443            // 478
        ,  1.861    ,  0.443            // 479
        ,  2.747    ,  1.329            // 480
        ,  2.569    ,  1.329            // 481
        ,  2.747    ,  1.152            // 482
        ,  2.569    ,  1.152            // 483
        ,  2.215    ,  1.329            // 484
        ,  2.392    ,  1.329            // 485
        ,  2.215    ,  1.152            // 486
        ,  2.392    ,  1.152            // 487
        ,  2.747    ,  0.797            // 488
        ,  2.569    ,  0.797            // 489
        ,  2.747    ,  0.975            // 490
        ,  2.569    ,  0.975            // 491
        ,  2.215    ,  0.797            // 492
        ,  2.392    ,  0.797            // 493
        ,  2.215    ,  0.975            // 494
        ,  2.392    ,  0.975            // 495
        ,  1.506    ,  1.329            // 496
        ,  1.683    ,  1.329            // 497
        ,  1.506    ,  1.152            // 498
        ,  1.683    ,  1.152            // 499
        ,  2.038    ,  1.329            // 500
        ,  1.861    ,  1.329            // 501
        ,  2.038    ,  1.152            // 502
        ,  1.861    ,  1.152            // 503
        ,  1.506    ,  0.797            // 504
        ,  1.683    ,  0.797            // 505
        ,  1.506    ,  0.975            // 506
        ,  1.683    ,  0.975            // 507
        ,  2.038    ,  0.797            // 508
        ,  1.861    ,  0.797            // 509
        ,  2.038    ,  0.975            // 510
        ,  1.861    ,  0.975            // 511
        ,  2.747    , -2.924            // 512
        ,  2.569    , -2.924            // 513
        ,  2.747    , -3.101            // 514
        ,  2.569    , -3.101            // 515
        ,  2.215    , -2.924            // 516
        ,  2.392    , -2.924            // 517
        ,  2.215    , -3.101            // 518
        ,  2.392    , -3.101            // 519
        ,  2.747    , -3.455            // 520
        ,  2.569    , -3.455            // 521
        ,  2.747    , -3.278            // 522
        ,  2.569    , -3.278            // 523
        ,  2.215    , -3.455            // 524
        ,  2.392    , -3.455            // 525
        ,  2.215    , -3.278            // 526
        ,  2.392    , -3.278            // 527
        ,  1.506    , -2.924            // 528
        ,  1.683    , -2.924            // 529
        ,  1.506    , -3.101            // 530
        ,  1.683    , -3.101            // 531
        ,  2.038    , -2.924            // 532
        ,  1.861    , -2.924            // 533
        ,  2.038    , -3.101            // 534
        ,  1.861    , -3.101            // 535
        ,  1.506    , -3.455            // 536
        ,  1.683    , -3.455            // 537
        ,  1.506    , -3.278            // 538
        ,  1.683    , -3.278            // 539
        ,  2.038    , -3.455            // 540
        ,  1.861    , -3.455            // 541
        ,  2.038    , -3.278            // 542
        ,  1.861    , -3.278            // 543
        ,  2.747    , -4.164            // 544
        ,  2.569    , -4.164            // 545
        ,  2.747    , -3.987            // 546
        ,  2.569    , -3.987            // 547
        ,  2.215    , -4.164            // 548
        ,  2.392    , -4.164            // 549
        ,  2.215    , -3.987            // 550
        ,  2.392    , -3.987            // 551
        ,  2.747    , -3.633            // 552
        ,  2.569    , -3.633            // 553
        ,  2.747    ,  -3.81            // 554
        ,  2.569    ,  -3.81            // 555
        ,  2.215    , -3.633            // 556
        ,  2.392    , -3.633            // 557
        ,  2.215    ,  -3.81            // 558
        ,  2.392    ,  -3.81            // 559
        ,  1.506    , -4.164            // 560
        ,  1.683    , -4.164            // 561
        ,  1.506    , -3.987            // 562
        ,  1.683    , -3.987            // 563
        ,  2.038    , -4.164            // 564
        ,  1.861    , -4.164            // 565
        ,  2.038    , -3.987            // 566
        ,  1.861    , -3.987            // 567
        ,  1.506    , -3.633            // 568
        ,  1.683    , -3.633            // 569
        ,  1.506    ,  -3.81            // 570
        ,  1.683    ,  -3.81            // 571
        ,  2.038    , -3.633            // 572
        ,  1.861    , -3.633            // 573
        ,  2.038    ,  -3.81            // 574
        ,  1.861    ,  -3.81            // 575
        ,  2.924    , -2.747            // 576
        ,  3.101    , -2.747            // 577
        ,  2.924    , -2.569            // 578
        ,  3.101    , -2.569            // 579
        ,  3.455    , -2.747            // 580
        ,  3.278    , -2.747            // 581
        ,  3.455    , -2.569            // 582
        ,  3.278    , -2.569            // 583
        ,  2.924    , -2.215            // 584
        ,  3.101    , -2.215            // 585
        ,  2.924    , -2.392            // 586
        ,  3.101    , -2.392            // 587
        ,  3.455    , -2.215            // 588
        ,  3.278    , -2.215            // 589
        ,  3.455    , -2.392            // 590
        ,  3.278    , -2.392            // 591
        ,  4.164    , -2.747            // 592
        ,  3.987    , -2.747            // 593
        ,  4.164    , -2.569            // 594
        ,  3.987    , -2.569            // 595
        ,  3.633    , -2.747            // 596
        ,   3.81    , -2.747            // 597
        ,  3.633    , -2.569            // 598
        ,   3.81    , -2.569            // 599
        ,  4.164    , -2.215            // 600
        ,  3.987    , -2.215            // 601
        ,  4.164    , -2.392            // 602
        ,  3.987    , -2.392            // 603
        ,  3.633    , -2.215            // 604
        ,   3.81    , -2.215            // 605
        ,  3.633    , -2.392            // 606
        ,   3.81    , -2.392            // 607
        ,  2.924    , -1.506            // 608
        ,  3.101    , -1.506            // 609
        ,  2.924    , -1.683            // 610
        ,  3.101    , -1.683            // 611
        ,  3.455    , -1.506            // 612
        ,  3.278    , -1.506            // 613
        ,  3.455    , -1.683            // 614
        ,  3.278    , -1.683            // 615
        ,  2.924    , -2.038            // 616
        ,  3.101    , -2.038            // 617
        ,  2.924    , -1.861            // 618
        ,  3.101    , -1.861            // 619
        ,  3.455    , -2.038            // 620
        ,  3.278    , -2.038            // 621
        ,  3.455    , -1.861            // 622
        ,  3.278    , -1.861            // 623
        ,  4.164    , -1.506            // 624
        ,  3.987    , -1.506            // 625
        ,  4.164    , -1.683            // 626
        ,  3.987    , -1.683            // 627
        ,  3.633    , -1.506            // 628
        ,   3.81    , -1.506            // 629
        ,  3.633    , -1.683            // 630
        ,   3.81    , -1.683            // 631
        ,  4.164    , -2.038            // 632
        ,  3.987    , -2.038            // 633
        ,  4.164    , -1.861            // 634
        ,  3.987    , -1.861            // 635
        ,  3.633    , -2.038            // 636
        ,   3.81    , -2.038            // 637
        ,  3.633    , -1.861            // 638
        ,   3.81    , -1.861            // 639
        ,  0.089    , -2.924            // 640
        ,  0.266    , -2.924            // 641
        ,  0.089    , -3.101            // 642
        ,  0.266    , -3.101            // 643
        ,   0.62    , -2.924            // 644
        ,  0.443    , -2.924            // 645
        ,   0.62    , -3.101            // 646
        ,  0.443    , -3.101            // 647
        ,  0.089    , -3.455            // 648
        ,  0.266    , -3.455            // 649
        ,  0.089    , -3.278            // 650
        ,  0.266    , -3.278            // 651
        ,   0.62    , -3.455            // 652
        ,  0.443    , -3.455            // 653
        ,   0.62    , -3.278            // 654
        ,  0.443    , -3.278            // 655
        ,  1.329    , -2.924            // 656
        ,  1.152    , -2.924            // 657
        ,  1.329    , -3.101            // 658
        ,  1.152    , -3.101            // 659
        ,  0.797    , -2.924            // 660
        ,  0.975    , -2.924            // 661
        ,  0.797    , -3.101            // 662
        ,  0.975    , -3.101            // 663
        ,  1.329    , -3.455            // 664
        ,  1.152    , -3.455            // 665
        ,  1.329    , -3.278            // 666
        ,  1.152    , -3.278            // 667
        ,  0.797    , -3.455            // 668
        ,  0.975    , -3.455            // 669
        ,  0.797    , -3.278            // 670
        ,  0.975    , -3.278            // 671
        ,  0.089    , -4.164            // 672
        ,  0.266    , -4.164            // 673
        ,  0.089    , -3.987            // 674
        ,  0.266    , -3.987            // 675
        ,   0.62    , -4.164            // 676
        ,  0.443    , -4.164            // 677
        ,   0.62    , -3.987            // 678
        ,  0.443    , -3.987            // 679
        ,  0.089    , -3.633            // 680
        ,  0.266    , -3.633            // 681
        ,  0.089    ,  -3.81            // 682
        ,  0.266    ,  -3.81            // 683
        ,   0.62    , -3.633            // 684
        ,  0.443    , -3.633            // 685
        ,   0.62    ,  -3.81            // 686
        ,  0.443    ,  -3.81            // 687
        ,  1.329    , -4.164            // 688
        ,  1.152    , -4.164            // 689
        ,  1.329    , -3.987            // 690
        ,  1.152    , -3.987            // 691
        ,  0.797    , -4.164            // 692
        ,  0.975    , -4.164            // 693
        ,  0.797    , -3.987            // 694
        ,  0.975    , -3.987            // 695
        ,  1.329    , -3.633            // 696
        ,  1.152    , -3.633            // 697
        ,  1.329    ,  -3.81            // 698
        ,  1.152    ,  -3.81            // 699
        ,  0.797    , -3.633            // 700
        ,  0.975    , -3.633            // 701
        ,  0.797    ,  -3.81            // 702
        ,  0.975    ,  -3.81            // 703
        ,  2.924    , -0.089            // 704
        ,  3.101    , -0.089            // 705
        ,  2.924    , -0.266            // 706
        ,  3.101    , -0.266            // 707
        ,  3.455    , -0.089            // 708
        ,  3.278    , -0.089            // 709
        ,  3.455    , -0.266            // 710
        ,  3.278    , -0.266            // 711
        ,  2.924    ,  -0.62            // 712
        ,  3.101    ,  -0.62            // 713
        ,  2.924    , -0.443            // 714
        ,  3.101    , -0.443            // 715
        ,  3.455    ,  -0.62            // 716
        ,  3.278    ,  -0.62            // 717
        ,  3.455    , -0.443            // 718
        ,  3.278    , -0.443            // 719
        ,  4.164    , -0.089            // 720
        ,  3.987    , -0.089            // 721
        ,  4.164    , -0.266            // 722
        ,  3.987    , -0.266            // 723
        ,  3.633    , -0.089            // 724
        ,   3.81    , -0.089            // 725
        ,  3.633    , -0.266            // 726
        ,   3.81    , -0.266            // 727
        ,  4.164    ,  -0.62            // 728
        ,  3.987    ,  -0.62            // 729
        ,  4.164    , -0.443            // 730
        ,  3.987    , -0.443            // 731
        ,  3.633    ,  -0.62            // 732
        ,   3.81    ,  -0.62            // 733
        ,  3.633    , -0.443            // 734
        ,   3.81    , -0.443            // 735
        ,  2.924    , -1.329            // 736
        ,  3.101    , -1.329            // 737
        ,  2.924    , -1.152            // 738
        ,  3.101    , -1.152            // 739
        ,  3.455    , -1.329            // 740
        ,  3.278    , -1.329            // 741
        ,  3.455    , -1.152            // 742
        ,  3.278    , -1.152            // 743
        ,  2.924    , -0.797            // 744
        ,  3.101    , -0.797            // 745
        ,  2.924    , -0.975            // 746
        ,  3.101    , -0.975            // 747
        ,  3.455    , -0.797            // 748
        ,  3.278    , -0.797            // 749
        ,  3.455    , -0.975            // 750
        ,  3.278    , -0.975            // 751
        ,  4.164    , -1.329            // 752
        ,  3.987    , -1.329            // 753
        ,  4.164    , -1.152            // 754
        ,  3.987    , -1.152            // 755
        ,  3.633    , -1.329            // 756
        ,   3.81    , -1.329            // 757
        ,  3.633    , -1.152            // 758
        ,   3.81    , -1.152            // 759
        ,  4.164    , -0.797            // 760
        ,  3.987    , -0.797            // 761
        ,  4.164    , -0.975            // 762
        ,  3.987    , -0.975            // 763
        ,  3.633    , -0.797            // 764
        ,   3.81    , -0.797            // 765
        ,  3.633    , -0.975            // 766
        ,   3.81    , -0.975            // 767
        ,  0.089    , -2.747            // 768
        ,  0.266    , -2.747            // 769
        ,  0.089    , -2.569            // 770
        ,  0.266    , -2.569            // 771
        ,   0.62    , -2.747            // 772
        ,  0.443    , -2.747            // 773
        ,   0.62    , -2.569            // 774
        ,  0.443    , -2.569            // 775
        ,  0.089    , -2.215            // 776
        ,  0.266    , -2.215            // 777
        ,  0.089    , -2.392            // 778
        ,  0.266    , -2.392            // 779
        ,   0.62    , -2.215            // 780
        ,  0.443    , -2.215            // 781
        ,   0.62    , -2.392            // 782
        ,  0.443    , -2.392            // 783
        ,  1.329    , -2.747            // 784
        ,  1.152    , -2.747            // 785
        ,  1.329    , -2.569            // 786
        ,  1.152    , -2.569            // 787
        ,  0.797    , -2.747            // 788
        ,  0.975    , -2.747            // 789
        ,  0.797    , -2.569            // 790
        ,  0.975    , -2.569            // 791
        ,  1.329    , -2.215            // 792
        ,  1.152    , -2.215            // 793
        ,  1.329    , -2.392            // 794
        ,  1.152    , -2.392            // 795
        ,  0.797    , -2.215            // 796
        ,  0.975    , -2.215            // 797
        ,  0.797    , -2.392            // 798
        ,  0.975    , -2.392            // 799
        ,  0.089    , -1.506            // 800
        ,  0.266    , -1.506            // 801
        ,  0.089    , -1.683            // 802
        ,  0.266    , -1.683            // 803
        ,   0.62    , -1.506            // 804
        ,  0.443    , -1.506            // 805
        ,   0.62    , -1.683            // 806
        ,  0.443    , -1.683            // 807
        ,  0.089    , -2.038            // 808
        ,  0.266    , -2.038            // 809
        ,  0.089    , -1.861            // 810
        ,  0.266    , -1.861            // 811
        ,   0.62    , -2.038            // 812
        ,  0.443    , -2.038            // 813
        ,   0.62    , -1.861            // 814
        ,  0.443    , -1.861            // 815
        ,  1.329    , -1.506            // 816
        ,  1.152    , -1.506            // 817
        ,  1.329    , -1.683            // 818
        ,  1.152    , -1.683            // 819
        ,  0.797    , -1.506            // 820
        ,  0.975    , -1.506            // 821
        ,  0.797    , -1.683            // 822
        ,  0.975    , -1.683            // 823
        ,  1.329    , -2.038            // 824
        ,  1.152    , -2.038            // 825
        ,  1.329    , -1.861            // 826
        ,  1.152    , -1.861            // 827
        ,  0.797    , -2.038            // 828
        ,  0.975    , -2.038            // 829
        ,  0.797    , -1.861            // 830
        ,  0.975    , -1.861            // 831
        ,  2.747    , -2.747            // 832
        ,  2.569    , -2.747            // 833
        ,  2.747    , -2.569            // 834
        ,  2.569    , -2.569            // 835
        ,  2.215    , -2.747            // 836
        ,  2.392    , -2.747            // 837
        ,  2.215    , -2.569            // 838
        ,  2.392    , -2.569            // 839
        ,  2.747    , -2.215            // 840
        ,  2.569    , -2.215            // 841
        ,  2.747    , -2.392            // 842
        ,  2.569    , -2.392            // 843
        ,  2.215    , -2.215            // 844
        ,  2.392    , -2.215            // 845
        ,  2.215    , -2.392            // 846
        ,  2.392    , -2.392            // 847
        ,  1.506    , -2.747            // 848
        ,  1.683    , -2.747            // 849
        ,  1.506    , -2.569            // 850
        ,  1.683    , -2.569            // 851
        ,  2.038    , -2.747            // 852
        ,  1.861    , -2.747            // 853
        ,  2.038    , -2.569            // 854
        ,  1.861    , -2.569            // 855
        ,  1.506    , -2.215            // 856
        ,  1.683    , -2.215            // 857
        ,  1.506    , -2.392            // 858
        ,  1.683    , -2.392            // 859
        ,  2.038    , -2.215            // 860
        ,  1.861    , -2.215            // 861
        ,  2.038    , -2.392            // 862
        ,  1.861    , -2.392            // 863
        ,  2.747    , -1.506            // 864
        ,  2.569    , -1.506            // 865
        ,  2.747    , -1.683            // 866
        ,  2.569    , -1.683            // 867
        ,  2.215    , -1.506            // 868
        ,  2.392    , -1.506            // 869
        ,  2.215    , -1.683            // 870
        ,  2.392    , -1.683            // 871
        ,  2.747    , -2.038            // 872
        ,  2.569    , -2.038            // 873
        ,  2.747    , -1.861            // 874
        ,  2.569    , -1.861            // 875
        ,  2.215    , -2.038            // 876
        ,  2.392    , -2.038            // 877
        ,  2.215    , -1.861            // 878
        ,  2.392    , -1.861            // 879
        ,  1.506    , -1.506            // 880
        ,  1.683    , -1.506            // 881
        ,  1.506    , -1.683            // 882
        ,  1.683    , -1.683            // 883
        ,  2.038    , -1.506            // 884
        ,  1.861    , -1.506            // 885
        ,  2.038    , -1.683            // 886
        ,  1.861    , -1.683            // 887
        ,  1.506    , -2.038            // 888
        ,  1.683    , -2.038            // 889
        ,  1.506    , -1.861            // 890
        ,  1.683    , -1.861            // 891
        ,  2.038    , -2.038            // 892
        ,  1.861    , -2.038            // 893
        ,  2.038    , -1.861            // 894
        ,  1.861    , -1.861            // 895
        ,  0.089    , -0.089            // 896
        ,  0.266    , -0.089            // 897
        ,  0.089    , -0.266            // 898
        ,  0.266    , -0.266            // 899
        ,   0.62    , -0.089            // 900
        ,  0.443    , -0.089            // 901
        ,   0.62    , -0.266            // 902
        ,  0.443    , -0.266            // 903
        ,  0.089    ,  -0.62            // 904
        ,  0.266    ,  -0.62            // 905
        ,  0.089    , -0.443            // 906
        ,  0.266    , -0.443            // 907
        ,   0.62    ,  -0.62            // 908
        ,  0.443    ,  -0.62            // 909
        ,   0.62    , -0.443            // 910
        ,  0.443    , -0.443            // 911
        ,  1.329    , -0.089            // 912
        ,  1.152    , -0.089            // 913
        ,  1.329    , -0.266            // 914
        ,  1.152    , -0.266            // 915
        ,  0.797    , -0.089            // 916
        ,  0.975    , -0.089            // 917
        ,  0.797    , -0.266            // 918
        ,  0.975    , -0.266            // 919
        ,  1.329    ,  -0.62            // 920
        ,  1.152    ,  -0.62            // 921
        ,  1.329    , -0.443            // 922
        ,  1.152    , -0.443            // 923
        ,  0.797    ,  -0.62            // 924
        ,  0.975    ,  -0.62            // 925
        ,  0.797    , -0.443            // 926
        ,  0.975    , -0.443            // 927
        ,  0.089    , -1.329            // 928
        ,  0.266    , -1.329            // 929
        ,  0.089    , -1.152            // 930
        ,  0.266    , -1.152            // 931
        ,   0.62    , -1.329            // 932
        ,  0.443    , -1.329            // 933
        ,   0.62    , -1.152            // 934
        ,  0.443    , -1.152            // 935
        ,  0.089    , -0.797            // 936
        ,  0.266    , -0.797            // 937
        ,  0.089    , -0.975            // 938
        ,  0.266    , -0.975            // 939
        ,   0.62    , -0.797            // 940
        ,  0.443    , -0.797            // 941
        ,   0.62    , -0.975            // 942
        ,  0.443    , -0.975            // 943
        ,  1.329    , -1.329            // 944
        ,  1.152    , -1.329            // 945
        ,  1.329    , -1.152            // 946
        ,  1.152    , -1.152            // 947
        ,  0.797    , -1.329            // 948
        ,  0.975    , -1.329            // 949
        ,  0.797    , -1.152            // 950
        ,  0.975    , -1.152            // 951
        ,  1.329    , -0.797            // 952
        ,  1.152    , -0.797            // 953
        ,  1.329    , -0.975            // 954
        ,  1.152    , -0.975            // 955
        ,  0.797    , -0.797            // 956
        ,  0.975    , -0.797            // 957
        ,  0.797    , -0.975            // 958
        ,  0.975    , -0.975            // 959
        ,  2.747    , -0.089            // 960
        ,  2.569    , -0.089            // 961
        ,  2.747    , -0.266            // 962
        ,  2.569    , -0.266            // 963
        ,  2.215    , -0.089            // 964
        ,  2.392    , -0.089            // 965
        ,  2.215    , -0.266            // 966
        ,  2.392    , -0.266            // 967
        ,  2.747    ,  -0.62            // 968
        ,  2.569    ,  -0.62            // 969
        ,  2.747    , -0.443            // 970
        ,  2.569    , -0.443            // 971
        ,  2.215    ,  -0.62            // 972
        ,  2.392    ,  -0.62            // 973
        ,  2.215    , -0.443            // 974
        ,  2.392    , -0.443            // 975
        ,  1.506    , -0.089            // 976
        ,  1.683    , -0.089            // 977
        ,  1.506    , -0.266            // 978
        ,  1.683    , -0.266            // 979
        ,  2.038    , -0.089            // 980
        ,  1.861    , -0.089            // 981
        ,  2.038    , -0.266            // 982
        ,  1.861    , -0.266            // 983
        ,  1.506    ,  -0.62            // 984
        ,  1.683    ,  -0.62            // 985
        ,  1.506    , -0.443            // 986
        ,  1.683    , -0.443            // 987
        ,  2.038    ,  -0.62            // 988
        ,  1.861    ,  -0.62            // 989
        ,  2.038    , -0.443            // 990
        ,  1.861    , -0.443            // 991
        ,  2.747    , -1.329            // 992
        ,  2.569    , -1.329            // 993
        ,  2.747    , -1.152            // 994
        ,  2.569    , -1.152            // 995
        ,  2.215    , -1.329            // 996
        ,  2.392    , -1.329            // 997
        ,  2.215    , -1.152            // 998
        ,  2.392    , -1.152            // 999
        ,  2.747    , -0.797            // 1000
        ,  2.569    , -0.797            // 1001
        ,  2.747    , -0.975            // 1002
        ,  2.569    , -0.975            // 1003
        ,  2.215    , -0.797            // 1004
        ,  2.392    , -0.797            // 1005
        ,  2.215    , -0.975            // 1006
        ,  2.392    , -0.975            // 1007
        ,  1.506    , -1.329            // 1008
        ,  1.683    , -1.329            // 1009
        ,  1.506    , -1.152            // 1010
        ,  1.683    , -1.152            // 1011
        ,  2.038    , -1.329            // 1012
        ,  1.861    , -1.329            // 1013
        ,  2.038    , -1.152            // 1014
        ,  1.861    , -1.152            // 1015
        ,  1.506    , -0.797            // 1016
        ,  1.683    , -0.797            // 1017
        ,  1.506    , -0.975            // 1018
        ,  1.683    , -0.975            // 1019
        ,  2.038    , -0.797            // 1020
        ,  1.861    , -0.797            // 1021
        ,  2.038    , -0.975            // 1022
        ,  1.861    , -0.975            // 1023
        , -2.747    ,  2.924            // 1024
        , -2.569    ,  2.924            // 1025
        , -2.747    ,  3.101            // 1026
        , -2.569    ,  3.101            // 1027
        , -2.215    ,  2.924            // 1028
        , -2.392    ,  2.924            // 1029
        , -2.215    ,  3.101            // 1030
        , -2.392    ,  3.101            // 1031
        , -2.747    ,  3.455            // 1032
        , -2.569    ,  3.455            // 1033
        , -2.747    ,  3.278            // 1034
        , -2.569    ,  3.278            // 1035
        , -2.215    ,  3.455            // 1036
        , -2.392    ,  3.455            // 1037
        , -2.215    ,  3.278            // 1038
        , -2.392    ,  3.278            // 1039
        , -1.506    ,  2.924            // 1040
        , -1.683    ,  2.924            // 1041
        , -1.506    ,  3.101            // 1042
        , -1.683    ,  3.101            // 1043
        , -2.038    ,  2.924            // 1044
        , -1.861    ,  2.924            // 1045
        , -2.038    ,  3.101            // 1046
        , -1.861    ,  3.101            // 1047
        , -1.506    ,  3.455            // 1048
        , -1.683    ,  3.455            // 1049
        , -1.506    ,  3.278            // 1050
        , -1.683    ,  3.278            // 1051
        , -2.038    ,  3.455            // 1052
        , -1.861    ,  3.455            // 1053
        , -2.038    ,  3.278            // 1054
        , -1.861    ,  3.278            // 1055
        , -2.747    ,  4.164            // 1056
        , -2.569    ,  4.164            // 1057
        , -2.747    ,  3.987            // 1058
        , -2.569    ,  3.987            // 1059
        , -2.215    ,  4.164            // 1060
        , -2.392    ,  4.164            // 1061
        , -2.215    ,  3.987            // 1062
        , -2.392    ,  3.987            // 1063
        , -2.747    ,  3.633            // 1064
        , -2.569    ,  3.633            // 1065
        , -2.747    ,   3.81            // 1066
        , -2.569    ,   3.81            // 1067
        , -2.215    ,  3.633            // 1068
        , -2.392    ,  3.633            // 1069
        , -2.215    ,   3.81            // 1070
        , -2.392    ,   3.81            // 1071
        , -1.506    ,  4.164            // 1072
        , -1.683    ,  4.164            // 1073
        , -1.506    ,  3.987            // 1074
        , -1.683    ,  3.987            // 1075
        , -2.038    ,  4.164            // 1076
        , -1.861    ,  4.164            // 1077
        , -2.038    ,  3.987            // 1078
        , -1.861    ,  3.987            // 1079
        , -1.506    ,  3.633            // 1080
        , -1.683    ,  3.633            // 1081
        , -1.506    ,   3.81            // 1082
        , -1.683    ,   3.81            // 1083
        , -2.038    ,  3.633            // 1084
        , -1.861    ,  3.633            // 1085
        , -2.038    ,   3.81            // 1086
        , -1.861    ,   3.81            // 1087
        , -2.924    ,  2.747            // 1088
        , -3.101    ,  2.747            // 1089
        , -2.924    ,  2.569            // 1090
        , -3.101    ,  2.569            // 1091
        , -3.455    ,  2.747            // 1092
        , -3.278    ,  2.747            // 1093
        , -3.455    ,  2.569            // 1094
        , -3.278    ,  2.569            // 1095
        , -2.924    ,  2.215            // 1096
        , -3.101    ,  2.215            // 1097
        , -2.924    ,  2.392            // 1098
        , -3.101    ,  2.392            // 1099
        , -3.455    ,  2.215            // 1100
        , -3.278    ,  2.215            // 1101
        , -3.455    ,  2.392            // 1102
        , -3.278    ,  2.392            // 1103
        , -4.164    ,  2.747            // 1104
        , -3.987    ,  2.747            // 1105
        , -4.164    ,  2.569            // 1106
        , -3.987    ,  2.569            // 1107
        , -3.633    ,  2.747            // 1108
        ,  -3.81    ,  2.747            // 1109
        , -3.633    ,  2.569            // 1110
        ,  -3.81    ,  2.569            // 1111
        , -4.164    ,  2.215            // 1112
        , -3.987    ,  2.215            // 1113
        , -4.164    ,  2.392            // 1114
        , -3.987    ,  2.392            // 1115
        , -3.633    ,  2.215            // 1116
        ,  -3.81    ,  2.215            // 1117
        , -3.633    ,  2.392            // 1118
        ,  -3.81    ,  2.392            // 1119
        , -2.924    ,  1.506            // 1120
        , -3.101    ,  1.506            // 1121
        , -2.924    ,  1.683            // 1122
        , -3.101    ,  1.683            // 1123
        , -3.455    ,  1.506            // 1124
        , -3.278    ,  1.506            // 1125
        , -3.455    ,  1.683            // 1126
        , -3.278    ,  1.683            // 1127
        , -2.924    ,  2.038            // 1128
        , -3.101    ,  2.038            // 1129
        , -2.924    ,  1.861            // 1130
        , -3.101    ,  1.861            // 1131
        , -3.455    ,  2.038            // 1132
        , -3.278    ,  2.038            // 1133
        , -3.455    ,  1.861            // 1134
        , -3.278    ,  1.861            // 1135
        , -4.164    ,  1.506            // 1136
        , -3.987    ,  1.506            // 1137
        , -4.164    ,  1.683            // 1138
        , -3.987    ,  1.683            // 1139
        , -3.633    ,  1.506            // 1140
        ,  -3.81    ,  1.506            // 1141
        , -3.633    ,  1.683            // 1142
        ,  -3.81    ,  1.683            // 1143
        , -4.164    ,  2.038            // 1144
        , -3.987    ,  2.038            // 1145
        , -4.164    ,  1.861            // 1146
        , -3.987    ,  1.861            // 1147
        , -3.633    ,  2.038            // 1148
        ,  -3.81    ,  2.038            // 1149
        , -3.633    ,  1.861            // 1150
        ,  -3.81    ,  1.861            // 1151
        , -0.089    ,  2.924            // 1152
        , -0.266    ,  2.924            // 1153
        , -0.089    ,  3.101            // 1154
        , -0.266    ,  3.101            // 1155
        ,  -0.62    ,  2.924            // 1156
        , -0.443    ,  2.924            // 1157
        ,  -0.62    ,  3.101            // 1158
        , -0.443    ,  3.101            // 1159
        , -0.089    ,  3.455            // 1160
        , -0.266    ,  3.455            // 1161
        , -0.089    ,  3.278            // 1162
        , -0.266    ,  3.278            // 1163
        ,  -0.62    ,  3.455            // 1164
        , -0.443    ,  3.455            // 1165
        ,  -0.62    ,  3.278            // 1166
        , -0.443    ,  3.278            // 1167
        , -1.329    ,  2.924            // 1168
        , -1.152    ,  2.924            // 1169
        , -1.329    ,  3.101            // 1170
        , -1.152    ,  3.101            // 1171
        , -0.797    ,  2.924            // 1172
        , -0.975    ,  2.924            // 1173
        , -0.797    ,  3.101            // 1174
        , -0.975    ,  3.101            // 1175
        , -1.329    ,  3.455            // 1176
        , -1.152    ,  3.455            // 1177
        , -1.329    ,  3.278            // 1178
        , -1.152    ,  3.278            // 1179
        , -0.797    ,  3.455            // 1180
        , -0.975    ,  3.455            // 1181
        , -0.797    ,  3.278            // 1182
        , -0.975    ,  3.278            // 1183
        , -0.089    ,  4.164            // 1184
        , -0.266    ,  4.164            // 1185
        , -0.089    ,  3.987            // 1186
        , -0.266    ,  3.987            // 1187
        ,  -0.62    ,  4.164            // 1188
        , -0.443    ,  4.164            // 1189
        ,  -0.62    ,  3.987            // 1190
        , -0.443    ,  3.987            // 1191
        , -0.089    ,  3.633            // 1192
        , -0.266    ,  3.633            // 1193
        , -0.089    ,   3.81            // 1194
        , -0.266    ,   3.81            // 1195
        ,  -0.62    ,  3.633            // 1196
        , -0.443    ,  3.633            // 1197
        ,  -0.62    ,   3.81            // 1198
        , -0.443    ,   3.81            // 1199
        , -1.329    ,  4.164            // 1200
        , -1.152    ,  4.164            // 1201
        , -1.329    ,  3.987            // 1202
        , -1.152    ,  3.987            // 1203
        , -0.797    ,  4.164            // 1204
        , -0.975    ,  4.164            // 1205
        , -0.797    ,  3.987            // 1206
        , -0.975    ,  3.987            // 1207
        , -1.329    ,  3.633            // 1208
        , -1.152    ,  3.633            // 1209
        , -1.329    ,   3.81            // 1210
        , -1.152    ,   3.81            // 1211
        , -0.797    ,  3.633            // 1212
        , -0.975    ,  3.633            // 1213
        , -0.797    ,   3.81            // 1214
        , -0.975    ,   3.81            // 1215
        , -2.924    ,  0.089            // 1216
        , -3.101    ,  0.089            // 1217
        , -2.924    ,  0.266            // 1218
        , -3.101    ,  0.266            // 1219
        , -3.455    ,  0.089            // 1220
        , -3.278    ,  0.089            // 1221
        , -3.455    ,  0.266            // 1222
        , -3.278    ,  0.266            // 1223
        , -2.924    ,   0.62            // 1224
        , -3.101    ,   0.62            // 1225
        , -2.924    ,  0.443            // 1226
        , -3.101    ,  0.443            // 1227
        , -3.455    ,   0.62            // 1228
        , -3.278    ,   0.62            // 1229
        , -3.455    ,  0.443            // 1230
        , -3.278    ,  0.443            // 1231
        , -4.164    ,  0.089            // 1232
        , -3.987    ,  0.089            // 1233
        , -4.164    ,  0.266            // 1234
        , -3.987    ,  0.266            // 1235
        , -3.633    ,  0.089            // 1236
        ,  -3.81    ,  0.089            // 1237
        , -3.633    ,  0.266            // 1238
        ,  -3.81    ,  0.266            // 1239
        , -4.164    ,   0.62            // 1240
        , -3.987    ,   0.62            // 1241
        , -4.164    ,  0.443            // 1242
        , -3.987    ,  0.443            // 1243
        , -3.633    ,   0.62            // 1244
        ,  -3.81    ,   0.62            // 1245
        , -3.633    ,  0.443            // 1246
        ,  -3.81    ,  0.443            // 1247
        , -2.924    ,  1.329            // 1248
        , -3.101    ,  1.329            // 1249
        , -2.924    ,  1.152            // 1250
        , -3.101    ,  1.152            // 1251
        , -3.455    ,  1.329            // 1252
        , -3.278    ,  1.329            // 1253
        , -3.455    ,  1.152            // 1254
        , -3.278    ,  1.152            // 1255
        , -2.924    ,  0.797            // 1256
        , -3.101    ,  0.797            // 1257
        , -2.924    ,  0.975            // 1258
        , -3.101    ,  0.975            // 1259
        , -3.455    ,  0.797            // 1260
        , -3.278    ,  0.797            // 1261
        , -3.455    ,  0.975            // 1262
        , -3.278    ,  0.975            // 1263
        , -4.164    ,  1.329            // 1264
        , -3.987    ,  1.329            // 1265
        , -4.164    ,  1.152            // 1266
        , -3.987    ,  1.152            // 1267
        , -3.633    ,  1.329            // 1268
        ,  -3.81    ,  1.329            // 1269
        , -3.633    ,  1.152            // 1270
        ,  -3.81    ,  1.152            // 1271
        , -4.164    ,  0.797            // 1272
        , -3.987    ,  0.797            // 1273
        , -4.164    ,  0.975            // 1274
        , -3.987    ,  0.975            // 1275
        , -3.633    ,  0.797            // 1276
        ,  -3.81    ,  0.797            // 1277
        , -3.633    ,  0.975            // 1278
        ,  -3.81    ,  0.975            // 1279
        , -0.089    ,  2.747            // 1280
        , -0.266    ,  2.747            // 1281
        , -0.089    ,  2.569            // 1282
        , -0.266    ,  2.569            // 1283
        ,  -0.62    ,  2.747            // 1284
        , -0.443    ,  2.747            // 1285
        ,  -0.62    ,  2.569            // 1286
        , -0.443    ,  2.569            // 1287
        , -0.089    ,  2.215            // 1288
        , -0.266    ,  2.215            // 1289
        , -0.089    ,  2.392            // 1290
        , -0.266    ,  2.392            // 1291
        ,  -0.62    ,  2.215            // 1292
        , -0.443    ,  2.215            // 1293
        ,  -0.62    ,  2.392            // 1294
        , -0.443    ,  2.392            // 1295
        , -1.329    ,  2.747            // 1296
        , -1.152    ,  2.747            // 1297
        , -1.329    ,  2.569            // 1298
        , -1.152    ,  2.569            // 1299
        , -0.797    ,  2.747            // 1300
        , -0.975    ,  2.747            // 1301
        , -0.797    ,  2.569            // 1302
        , -0.975    ,  2.569            // 1303
        , -1.329    ,  2.215            // 1304
        , -1.152    ,  2.215            // 1305
        , -1.329    ,  2.392            // 1306
        , -1.152    ,  2.392            // 1307
        , -0.797    ,  2.215            // 1308
        , -0.975    ,  2.215            // 1309
        , -0.797    ,  2.392            // 1310
        , -0.975    ,  2.392            // 1311
        , -0.089    ,  1.506            // 1312
        , -0.266    ,  1.506            // 1313
        , -0.089    ,  1.683            // 1314
        , -0.266    ,  1.683            // 1315
        ,  -0.62    ,  1.506            // 1316
        , -0.443    ,  1.506            // 1317
        ,  -0.62    ,  1.683            // 1318
        , -0.443    ,  1.683            // 1319
        , -0.089    ,  2.038            // 1320
        , -0.266    ,  2.038            // 1321
        , -0.089    ,  1.861            // 1322
        , -0.266    ,  1.861            // 1323
        ,  -0.62    ,  2.038            // 1324
        , -0.443    ,  2.038            // 1325
        ,  -0.62    ,  1.861            // 1326
        , -0.443    ,  1.861            // 1327
        , -1.329    ,  1.506            // 1328
        , -1.152    ,  1.506            // 1329
        , -1.329    ,  1.683            // 1330
        , -1.152    ,  1.683            // 1331
        , -0.797    ,  1.506            // 1332
        , -0.975    ,  1.506            // 1333
        , -0.797    ,  1.683            // 1334
        , -0.975    ,  1.683            // 1335
        , -1.329    ,  2.038            // 1336
        , -1.152    ,  2.038            // 1337
        , -1.329    ,  1.861            // 1338
        , -1.152    ,  1.861            // 1339
        , -0.797    ,  2.038            // 1340
        , -0.975    ,  2.038            // 1341
        , -0.797    ,  1.861            // 1342
        , -0.975    ,  1.861            // 1343
        , -2.747    ,  2.747            // 1344
        , -2.569    ,  2.747            // 1345
        , -2.747    ,  2.569            // 1346
        , -2.569    ,  2.569            // 1347
        , -2.215    ,  2.747            // 1348
        , -2.392    ,  2.747            // 1349
        , -2.215    ,  2.569            // 1350
        , -2.392    ,  2.569            // 1351
        , -2.747    ,  2.215            // 1352
        , -2.569    ,  2.215            // 1353
        , -2.747    ,  2.392            // 1354
        , -2.569    ,  2.392            // 1355
        , -2.215    ,  2.215            // 1356
        , -2.392    ,  2.215            // 1357
        , -2.215    ,  2.392            // 1358
        , -2.392    ,  2.392            // 1359
        , -1.506    ,  2.747            // 1360
        , -1.683    ,  2.747            // 1361
        , -1.506    ,  2.569            // 1362
        , -1.683    ,  2.569            // 1363
        , -2.038    ,  2.747            // 1364
        , -1.861    ,  2.747            // 1365
        , -2.038    ,  2.569            // 1366
        , -1.861    ,  2.569            // 1367
        , -1.506    ,  2.215            // 1368
        , -1.683    ,  2.215            // 1369
        , -1.506    ,  2.392            // 1370
        , -1.683    ,  2.392            // 1371
        , -2.038    ,  2.215            // 1372
        , -1.861    ,  2.215            // 1373
        , -2.038    ,  2.392            // 1374
        , -1.861    ,  2.392            // 1375
        , -2.747    ,  1.506            // 1376
        , -2.569    ,  1.506            // 1377
        , -2.747    ,  1.683            // 1378
        , -2.569    ,  1.683            // 1379
        , -2.215    ,  1.506            // 1380
        , -2.392    ,  1.506            // 1381
        , -2.215    ,  1.683            // 1382
        , -2.392    ,  1.683            // 1383
        , -2.747    ,  2.038            // 1384
        , -2.569    ,  2.038            // 1385
        , -2.747    ,  1.861            // 1386
        , -2.569    ,  1.861            // 1387
        , -2.215    ,  2.038            // 1388
        , -2.392    ,  2.038            // 1389
        , -2.215    ,  1.861            // 1390
        , -2.392    ,  1.861            // 1391
        , -1.506    ,  1.506            // 1392
        , -1.683    ,  1.506            // 1393
        , -1.506    ,  1.683            // 1394
        , -1.683    ,  1.683            // 1395
        , -2.038    ,  1.506            // 1396
        , -1.861    ,  1.506            // 1397
        , -2.038    ,  1.683            // 1398
        , -1.861    ,  1.683            // 1399
        , -1.506    ,  2.038            // 1400
        , -1.683    ,  2.038            // 1401
        , -1.506    ,  1.861            // 1402
        , -1.683    ,  1.861            // 1403
        , -2.038    ,  2.038            // 1404
        , -1.861    ,  2.038            // 1405
        , -2.038    ,  1.861            // 1406
        , -1.861    ,  1.861            // 1407
        , -0.089    ,  0.089            // 1408
        , -0.266    ,  0.089            // 1409
        , -0.089    ,  0.266            // 1410
        , -0.266    ,  0.266            // 1411
        ,  -0.62    ,  0.089            // 1412
        , -0.443    ,  0.089            // 1413
        ,  -0.62    ,  0.266            // 1414
        , -0.443    ,  0.266            // 1415
        , -0.089    ,   0.62            // 1416
        , -0.266    ,   0.62            // 1417
        , -0.089    ,  0.443            // 1418
        , -0.266    ,  0.443            // 1419
        ,  -0.62    ,   0.62            // 1420
        , -0.443    ,   0.62            // 1421
        ,  -0.62    ,  0.443            // 1422
        , -0.443    ,  0.443            // 1423
        , -1.329    ,  0.089            // 1424
        , -1.152    ,  0.089            // 1425
        , -1.329    ,  0.266            // 1426
        , -1.152    ,  0.266            // 1427
        , -0.797    ,  0.089            // 1428
        , -0.975    ,  0.089            // 1429
        , -0.797    ,  0.266            // 1430
        , -0.975    ,  0.266            // 1431
        , -1.329    ,   0.62            // 1432
        , -1.152    ,   0.62            // 1433
        , -1.329    ,  0.443            // 1434
        , -1.152    ,  0.443            // 1435
        , -0.797    ,   0.62            // 1436
        , -0.975    ,   0.62            // 1437
        , -0.797    ,  0.443            // 1438
        , -0.975    ,  0.443            // 1439
        , -0.089    ,  1.329            // 1440
        , -0.266    ,  1.329            // 1441
        , -0.089    ,  1.152            // 1442
        , -0.266    ,  1.152            // 1443
        ,  -0.62    ,  1.329            // 1444
        , -0.443    ,  1.329            // 1445
        ,  -0.62    ,  1.152            // 1446
        , -0.443    ,  1.152            // 1447
        , -0.089    ,  0.797            // 1448
        , -0.266    ,  0.797            // 1449
        , -0.089    ,  0.975            // 1450
        , -0.266    ,  0.975            // 1451
        ,  -0.62    ,  0.797            // 1452
        , -0.443    ,  0.797            // 1453
        ,  -0.62    ,  0.975            // 1454
        , -0.443    ,  0.975            // 1455
        , -1.329    ,  1.329            // 1456
        , -1.152    ,  1.329            // 1457
        , -1.329    ,  1.152            // 1458
        , -1.152    ,  1.152            // 1459
        , -0.797    ,  1.329            // 1460
        , -0.975    ,  1.329            // 1461
        , -0.797    ,  1.152            // 1462
        , -0.975    ,  1.152            // 1463
        , -1.329    ,  0.797            // 1464
        , -1.152    ,  0.797            // 1465
        , -1.329    ,  0.975            // 1466
        , -1.152    ,  0.975            // 1467
        , -0.797    ,  0.797            // 1468
        , -0.975    ,  0.797            // 1469
        , -0.797    ,  0.975            // 1470
        , -0.975    ,  0.975            // 1471
        , -2.747    ,  0.089            // 1472
        , -2.569    ,  0.089            // 1473
        , -2.747    ,  0.266            // 1474
        , -2.569    ,  0.266            // 1475
        , -2.215    ,  0.089            // 1476
        , -2.392    ,  0.089            // 1477
        , -2.215    ,  0.266            // 1478
        , -2.392    ,  0.266            // 1479
        , -2.747    ,   0.62            // 1480
        , -2.569    ,   0.62            // 1481
        , -2.747    ,  0.443            // 1482
        , -2.569    ,  0.443            // 1483
        , -2.215    ,   0.62            // 1484
        , -2.392    ,   0.62            // 1485
        , -2.215    ,  0.443            // 1486
        , -2.392    ,  0.443            // 1487
        , -1.506    ,  0.089            // 1488
        , -1.683    ,  0.089            // 1489
        , -1.506    ,  0.266            // 1490
        , -1.683    ,  0.266            // 1491
        , -2.038    ,  0.089            // 1492
        , -1.861    ,  0.089            // 1493
        , -2.038    ,  0.266            // 1494
        , -1.861    ,  0.266            // 1495
        , -1.506    ,   0.62            // 1496
        , -1.683    ,   0.62            // 1497
        , -1.506    ,  0.443            // 1498
        , -1.683    ,  0.443            // 1499
        , -2.038    ,   0.62            // 1500
        , -1.861    ,   0.62            // 1501
        , -2.038    ,  0.443            // 1502
        , -1.861    ,  0.443            // 1503
        , -2.747    ,  1.329            // 1504
        , -2.569    ,  1.329            // 1505
        , -2.747    ,  1.152            // 1506
        , -2.569    ,  1.152            // 1507
        , -2.215    ,  1.329            // 1508
        , -2.392    ,  1.329            // 1509
        , -2.215    ,  1.152            // 1510
        , -2.392    ,  1.152            // 1511
        , -2.747    ,  0.797            // 1512
        , -2.569    ,  0.797            // 1513
        , -2.747    ,  0.975            // 1514
        , -2.569    ,  0.975            // 1515
        , -2.215    ,  0.797            // 1516
        , -2.392    ,  0.797            // 1517
        , -2.215    ,  0.975            // 1518
        , -2.392    ,  0.975            // 1519
        , -1.506    ,  1.329            // 1520
        , -1.683    ,  1.329            // 1521
        , -1.506    ,  1.152            // 1522
        , -1.683    ,  1.152            // 1523
        , -2.038    ,  1.329            // 1524
        , -1.861    ,  1.329            // 1525
        , -2.038    ,  1.152            // 1526
        , -1.861    ,  1.152            // 1527
        , -1.506    ,  0.797            // 1528
        , -1.683    ,  0.797            // 1529
        , -1.506    ,  0.975            // 1530
        , -1.683    ,  0.975            // 1531
        , -2.038    ,  0.797            // 1532
        , -1.861    ,  0.797            // 1533
        , -2.038    ,  0.975            // 1534
        , -1.861    ,  0.975            // 1535
        , -2.747    , -2.924            // 1536
        , -2.569    , -2.924            // 1537
        , -2.747    , -3.101            // 1538
        , -2.569    , -3.101            // 1539
        , -2.215    , -2.924            // 1540
        , -2.392    , -2.924            // 1541
        , -2.215    , -3.101            // 1542
        , -2.392    , -3.101            // 1543
        , -2.747    , -3.455            // 1544
        , -2.569    , -3.455            // 1545
        , -2.747    , -3.278            // 1546
        , -2.569    , -3.278            // 1547
        , -2.215    , -3.455            // 1548
        , -2.392    , -3.455            // 1549
        , -2.215    , -3.278            // 1550
        , -2.392    , -3.278            // 1551
        , -1.506    , -2.924            // 1552
        , -1.683    , -2.924            // 1553
        , -1.506    , -3.101            // 1554
        , -1.683    , -3.101            // 1555
        , -2.038    , -2.924            // 1556
        , -1.861    , -2.924            // 1557
        , -2.038    , -3.101            // 1558
        , -1.861    , -3.101            // 1559
        , -1.506    , -3.455            // 1560
        , -1.683    , -3.455            // 1561
        , -1.506    , -3.278            // 1562
        , -1.683    , -3.278            // 1563
        , -2.038    , -3.455            // 1564
        , -1.861    , -3.455            // 1565
        , -2.038    , -3.278            // 1566
        , -1.861    , -3.278            // 1567
        , -2.747    , -4.164            // 1568
        , -2.569    , -4.164            // 1569
        , -2.747    , -3.987            // 1570
        , -2.569    , -3.987            // 1571
        , -2.215    , -4.164            // 1572
        , -2.392    , -4.164            // 1573
        , -2.215    , -3.987            // 1574
        , -2.392    , -3.987            // 1575
        , -2.747    , -3.633            // 1576
        , -2.569    , -3.633            // 1577
        , -2.747    ,  -3.81            // 1578
        , -2.569    ,  -3.81            // 1579
        , -2.215    , -3.633            // 1580
        , -2.392    , -3.633            // 1581
        , -2.215    ,  -3.81            // 1582
        , -2.392    ,  -3.81            // 1583
        , -1.506    , -4.164            // 1584
        , -1.683    , -4.164            // 1585
        , -1.506    , -3.987            // 1586
        , -1.683    , -3.987            // 1587
        , -2.038    , -4.164            // 1588
        , -1.861    , -4.164            // 1589
        , -2.038    , -3.987            // 1590
        , -1.861    , -3.987            // 1591
        , -1.506    , -3.633            // 1592
        , -1.683    , -3.633            // 1593
        , -1.506    ,  -3.81            // 1594
        , -1.683    ,  -3.81            // 1595
        , -2.038    , -3.633            // 1596
        , -1.861    , -3.633            // 1597
        , -2.038    ,  -3.81            // 1598
        , -1.861    ,  -3.81            // 1599
        , -2.924    , -2.747            // 1600
        , -3.101    , -2.747            // 1601
        , -2.924    , -2.569            // 1602
        , -3.101    , -2.569            // 1603
        , -3.455    , -2.747            // 1604
        , -3.278    , -2.747            // 1605
        , -3.455    , -2.569            // 1606
        , -3.278    , -2.569            // 1607
        , -2.924    , -2.215            // 1608
        , -3.101    , -2.215            // 1609
        , -2.924    , -2.392            // 1610
        , -3.101    , -2.392            // 1611
        , -3.455    , -2.215            // 1612
        , -3.278    , -2.215            // 1613
        , -3.455    , -2.392            // 1614
        , -3.278    , -2.392            // 1615
        , -4.164    , -2.747            // 1616
        , -3.987    , -2.747            // 1617
        , -4.164    , -2.569            // 1618
        , -3.987    , -2.569            // 1619
        , -3.633    , -2.747            // 1620
        ,  -3.81    , -2.747            // 1621
        , -3.633    , -2.569            // 1622
        ,  -3.81    , -2.569            // 1623
        , -4.164    , -2.215            // 1624
        , -3.987    , -2.215            // 1625
        , -4.164    , -2.392            // 1626
        , -3.987    , -2.392            // 1627
        , -3.633    , -2.215            // 1628
        ,  -3.81    , -2.215            // 1629
        , -3.633    , -2.392            // 1630
        ,  -3.81    , -2.392            // 1631
        , -2.924    , -1.506            // 1632
        , -3.101    , -1.506            // 1633
        , -2.924    , -1.683            // 1634
        , -3.101    , -1.683            // 1635
        , -3.455    , -1.506            // 1636
        , -3.278    , -1.506            // 1637
        , -3.455    , -1.683            // 1638
        , -3.278    , -1.683            // 1639
        , -2.924    , -2.038            // 1640
        , -3.101    , -2.038            // 1641
        , -2.924    , -1.861            // 1642
        , -3.101    , -1.861            // 1643
        , -3.455    , -2.038            // 1644
        , -3.278    , -2.038            // 1645
        , -3.455    , -1.861            // 1646
        , -3.278    , -1.861            // 1647
        , -4.164    , -1.506            // 1648
        , -3.987    , -1.506            // 1649
        , -4.164    , -1.683            // 1650
        , -3.987    , -1.683            // 1651
        , -3.633    , -1.506            // 1652
        ,  -3.81    , -1.506            // 1653
        , -3.633    , -1.683            // 1654
        ,  -3.81    , -1.683            // 1655
        , -4.164    , -2.038            // 1656
        , -3.987    , -2.038            // 1657
        , -4.164    , -1.861            // 1658
        , -3.987    , -1.861            // 1659
        , -3.633    , -2.038            // 1660
        ,  -3.81    , -2.038            // 1661
        , -3.633    , -1.861            // 1662
        ,  -3.81    , -1.861            // 1663
        , -0.089    , -2.924            // 1664
        , -0.266    , -2.924            // 1665
        , -0.089    , -3.101            // 1666
        , -0.266    , -3.101            // 1667
        ,  -0.62    , -2.924            // 1668
        , -0.443    , -2.924            // 1669
        ,  -0.62    , -3.101            // 1670
        , -0.443    , -3.101            // 1671
        , -0.089    , -3.455            // 1672
        , -0.266    , -3.455            // 1673
        , -0.089    , -3.278            // 1674
        , -0.266    , -3.278            // 1675
        ,  -0.62    , -3.455            // 1676
        , -0.443    , -3.455            // 1677
        ,  -0.62    , -3.278            // 1678
        , -0.443    , -3.278            // 1679
        , -1.329    , -2.924            // 1680
        , -1.152    , -2.924            // 1681
        , -1.329    , -3.101            // 1682
        , -1.152    , -3.101            // 1683
        , -0.797    , -2.924            // 1684
        , -0.975    , -2.924            // 1685
        , -0.797    , -3.101            // 1686
        , -0.975    , -3.101            // 1687
        , -1.329    , -3.455            // 1688
        , -1.152    , -3.455            // 1689
        , -1.329    , -3.278            // 1690
        , -1.152    , -3.278            // 1691
        , -0.797    , -3.455            // 1692
        , -0.975    , -3.455            // 1693
        , -0.797    , -3.278            // 1694
        , -0.975    , -3.278            // 1695
        , -0.089    , -4.164            // 1696
        , -0.266    , -4.164            // 1697
        , -0.089    , -3.987            // 1698
        , -0.266    , -3.987            // 1699
        ,  -0.62    , -4.164            // 1700
        , -0.443    , -4.164            // 1701
        ,  -0.62    , -3.987            // 1702
        , -0.443    , -3.987            // 1703
        , -0.089    , -3.633            // 1704
        , -0.266    , -3.633            // 1705
        , -0.089    ,  -3.81            // 1706
        , -0.266    ,  -3.81            // 1707
        ,  -0.62    , -3.633            // 1708
        , -0.443    , -3.633            // 1709
        ,  -0.62    ,  -3.81            // 1710
        , -0.443    ,  -3.81            // 1711
        , -1.329    , -4.164            // 1712
        , -1.152    , -4.164            // 1713
        , -1.329    , -3.987            // 1714
        , -1.152    , -3.987            // 1715
        , -0.797    , -4.164            // 1716
        , -0.975    , -4.164            // 1717
        , -0.797    , -3.987            // 1718
        , -0.975    , -3.987            // 1719
        , -1.329    , -3.633            // 1720
        , -1.152    , -3.633            // 1721
        , -1.329    ,  -3.81            // 1722
        , -1.152    ,  -3.81            // 1723
        , -0.797    , -3.633            // 1724
        , -0.975    , -3.633            // 1725
        , -0.797    ,  -3.81            // 1726
        , -0.975    ,  -3.81            // 1727
        , -2.924    , -0.089            // 1728
        , -3.101    , -0.089            // 1729
        , -2.924    , -0.266            // 1730
        , -3.101    , -0.266            // 1731
        , -3.455    , -0.089            // 1732
        , -3.278    , -0.089            // 1733
        , -3.455    , -0.266            // 1734
        , -3.278    , -0.266            // 1735
        , -2.924    ,  -0.62            // 1736
        , -3.101    ,  -0.62            // 1737
        , -2.924    , -0.443            // 1738
        , -3.101    , -0.443            // 1739
        , -3.455    ,  -0.62            // 1740
        , -3.278    ,  -0.62            // 1741
        , -3.455    , -0.443            // 1742
        , -3.278    , -0.443            // 1743
        , -4.164    , -0.089            // 1744
        , -3.987    , -0.089            // 1745
        , -4.164    , -0.266            // 1746
        , -3.987    , -0.266            // 1747
        , -3.633    , -0.089            // 1748
        ,  -3.81    , -0.089            // 1749
        , -3.633    , -0.266            // 1750
        ,  -3.81    , -0.266            // 1751
        , -4.164    ,  -0.62            // 1752
        , -3.987    ,  -0.62            // 1753
        , -4.164    , -0.443            // 1754
        , -3.987    , -0.443            // 1755
        , -3.633    ,  -0.62            // 1756
        ,  -3.81    ,  -0.62            // 1757
        , -3.633    , -0.443            // 1758
        ,  -3.81    , -0.443            // 1759
        , -2.924    , -1.329            // 1760
        , -3.101    , -1.329            // 1761
        , -2.924    , -1.152            // 1762
        , -3.101    , -1.152            // 1763
        , -3.455    , -1.329            // 1764
        , -3.278    , -1.329            // 1765
        , -3.455    , -1.152            // 1766
        , -3.278    , -1.152            // 1767
        , -2.924    , -0.797            // 1768
        , -3.101    , -0.797            // 1769
        , -2.924    , -0.975            // 1770
        , -3.101    , -0.975            // 1771
        , -3.455    , -0.797            // 1772
        , -3.278    , -0.797            // 1773
        , -3.455    , -0.975            // 1774
        , -3.278    , -0.975            // 1775
        , -4.164    , -1.329            // 1776
        , -3.987    , -1.329            // 1777
        , -4.164    , -1.152            // 1778
        , -3.987    , -1.152            // 1779
        , -3.633    , -1.329            // 1780
        ,  -3.81    , -1.329            // 1781
        , -3.633    , -1.152            // 1782
        ,  -3.81    , -1.152            // 1783
        , -4.164    , -0.797            // 1784
        , -3.987    , -0.797            // 1785
        , -4.164    , -0.975            // 1786
        , -3.987    , -0.975            // 1787
        , -3.633    , -0.797            // 1788
        ,  -3.81    , -0.797            // 1789
        , -3.633    , -0.975            // 1790
        ,  -3.81    , -0.975            // 1791
        , -0.089    , -2.747            // 1792
        , -0.266    , -2.747            // 1793
        , -0.089    , -2.569            // 1794
        , -0.266    , -2.569            // 1795
        ,  -0.62    , -2.747            // 1796
        , -0.443    , -2.747            // 1797
        ,  -0.62    , -2.569            // 1798
        , -0.443    , -2.569            // 1799
        , -0.089    , -2.215            // 1800
        , -0.266    , -2.215            // 1801
        , -0.089    , -2.392            // 1802
        , -0.266    , -2.392            // 1803
        ,  -0.62    , -2.215            // 1804
        , -0.443    , -2.215            // 1805
        ,  -0.62    , -2.392            // 1806
        , -0.443    , -2.392            // 1807
        , -1.329    , -2.747            // 1808
        , -1.152    , -2.747            // 1809
        , -1.329    , -2.569            // 1810
        , -1.152    , -2.569            // 1811
        , -0.797    , -2.747            // 1812
        , -0.975    , -2.747            // 1813
        , -0.797    , -2.569            // 1814
        , -0.975    , -2.569            // 1815
        , -1.329    , -2.215            // 1816
        , -1.152    , -2.215            // 1817
        , -1.329    , -2.392            // 1818
        , -1.152    , -2.392            // 1819
        , -0.797    , -2.215            // 1820
        , -0.975    , -2.215            // 1821
        , -0.797    , -2.392            // 1822
        , -0.975    , -2.392            // 1823
        , -0.089    , -1.506            // 1824
        , -0.266    , -1.506            // 1825
        , -0.089    , -1.683            // 1826
        , -0.266    , -1.683            // 1827
        ,  -0.62    , -1.506            // 1828
        , -0.443    , -1.506            // 1829
        ,  -0.62    , -1.683            // 1830
        , -0.443    , -1.683            // 1831
        , -0.089    , -2.038            // 1832
        , -0.266    , -2.038            // 1833
        , -0.089    , -1.861            // 1834
        , -0.266    , -1.861            // 1835
        ,  -0.62    , -2.038            // 1836
        , -0.443    , -2.038            // 1837
        ,  -0.62    , -1.861            // 1838
        , -0.443    , -1.861            // 1839
        , -1.329    , -1.506            // 1840
        , -1.152    , -1.506            // 1841
        , -1.329    , -1.683            // 1842
        , -1.152    , -1.683            // 1843
        , -0.797    , -1.506            // 1844
        , -0.975    , -1.506            // 1845
        , -0.797    , -1.683            // 1846
        , -0.975    , -1.683            // 1847
        , -1.329    , -2.038            // 1848
        , -1.152    , -2.038            // 1849
        , -1.329    , -1.861            // 1850
        , -1.152    , -1.861            // 1851
        , -0.797    , -2.038            // 1852
        , -0.975    , -2.038            // 1853
        , -0.797    , -1.861            // 1854
        , -0.975    , -1.861            // 1855
        , -2.747    , -2.747            // 1856
        , -2.569    , -2.747            // 1857
        , -2.747    , -2.569            // 1858
        , -2.569    , -2.569            // 1859
        , -2.215    , -2.747            // 1860
        , -2.392    , -2.747            // 1861
        , -2.215    , -2.569            // 1862
        , -2.392    , -2.569            // 1863
        , -2.747    , -2.215            // 1864
        , -2.569    , -2.215            // 1865
        , -2.747    , -2.392            // 1866
        , -2.569    , -2.392            // 1867
        , -2.215    , -2.215            // 1868
        , -2.392    , -2.215            // 1869
        , -2.215    , -2.392            // 1870
        , -2.392    , -2.392            // 1871
        , -1.506    , -2.747            // 1872
        , -1.683    , -2.747            // 1873
        , -1.506    , -2.569            // 1874
        , -1.683    , -2.569            // 1875
        , -2.038    , -2.747            // 1876
        , -1.861    , -2.747            // 1877
        , -2.038    , -2.569            // 1878
        , -1.861    , -2.569            // 1879
        , -1.506    , -2.215            // 1880
        , -1.683    , -2.215            // 1881
        , -1.506    , -2.392            // 1882
        , -1.683    , -2.392            // 1883
        , -2.038    , -2.215            // 1884
        , -1.861    , -2.215            // 1885
        , -2.038    , -2.392            // 1886
        , -1.861    , -2.392            // 1887
        , -2.747    , -1.506            // 1888
        , -2.569    , -1.506            // 1889
        , -2.747    , -1.683            // 1890
        , -2.569    , -1.683            // 1891
        , -2.215    , -1.506            // 1892
        , -2.392    , -1.506            // 1893
        , -2.215    , -1.683            // 1894
        , -2.392    , -1.683            // 1895
        , -2.747    , -2.038            // 1896
        , -2.569    , -2.038            // 1897
        , -2.747    , -1.861            // 1898
        , -2.569    , -1.861            // 1899
        , -2.215    , -2.038            // 1900
        , -2.392    , -2.038            // 1901
        , -2.215    , -1.861            // 1902
        , -2.392    , -1.861            // 1903
        , -1.506    , -1.506            // 1904
        , -1.683    , -1.506            // 1905
        , -1.506    , -1.683            // 1906
        , -1.683    , -1.683            // 1907
        , -2.038    , -1.506            // 1908
        , -1.861    , -1.506            // 1909
        , -2.038    , -1.683            // 1910
        , -1.861    , -1.683            // 1911
        , -1.506    , -2.038            // 1912
        , -1.683    , -2.038            // 1913
        , -1.506    , -1.861            // 1914
        , -1.683    , -1.861            // 1915
        , -2.038    , -2.038            // 1916
        , -1.861    , -2.038            // 1917
        , -2.038    , -1.861            // 1918
        , -1.861    , -1.861            // 1919
        , -0.089    , -0.089            // 1920
        , -0.266    , -0.089            // 1921
        , -0.089    , -0.266            // 1922
        , -0.266    , -0.266            // 1923
        ,  -0.62    , -0.089            // 1924
        , -0.443    , -0.089            // 1925
        ,  -0.62    , -0.266            // 1926
        , -0.443    , -0.266            // 1927
        , -0.089    ,  -0.62            // 1928
        , -0.266    ,  -0.62            // 1929
        , -0.089    , -0.443            // 1930
        , -0.266    , -0.443            // 1931
        ,  -0.62    ,  -0.62            // 1932
        , -0.443    ,  -0.62            // 1933
        ,  -0.62    , -0.443            // 1934
        , -0.443    , -0.443            // 1935
        , -1.329    , -0.089            // 1936
        , -1.152    , -0.089            // 1937
        , -1.329    , -0.266            // 1938
        , -1.152    , -0.266            // 1939
        , -0.797    , -0.089            // 1940
        , -0.975    , -0.089            // 1941
        , -0.797    , -0.266            // 1942
        , -0.975    , -0.266            // 1943
        , -1.329    ,  -0.62            // 1944
        , -1.152    ,  -0.62            // 1945
        , -1.329    , -0.443            // 1946
        , -1.152    , -0.443            // 1947
        , -0.797    ,  -0.62            // 1948
        , -0.975    ,  -0.62            // 1949
        , -0.797    , -0.443            // 1950
        , -0.975    , -0.443            // 1951
        , -0.089    , -1.329            // 1952
        , -0.266    , -1.329            // 1953
        , -0.089    , -1.152            // 1954
        , -0.266    , -1.152            // 1955
        ,  -0.62    , -1.329            // 1956
        , -0.443    , -1.329            // 1957
        ,  -0.62    , -1.152            // 1958
        , -0.443    , -1.152            // 1959
        , -0.089    , -0.797            // 1960
        , -0.266    , -0.797            // 1961
        , -0.089    , -0.975            // 1962
        , -0.266    , -0.975            // 1963
        ,  -0.62    , -0.797            // 1964
        , -0.443    , -0.797            // 1965
        ,  -0.62    , -0.975            // 1966
        , -0.443    , -0.975            // 1967
        , -1.329    , -1.329            // 1968
        , -1.152    , -1.329            // 1969
        , -1.329    , -1.152            // 1970
        , -1.152    , -1.152            // 1971
        , -0.797    , -1.329            // 1972
        , -0.975    , -1.329            // 1973
        , -0.797    , -1.152            // 1974
        , -0.975    , -1.152            // 1975
        , -1.329    , -0.797            // 1976
        , -1.152    , -0.797            // 1977
        , -1.329    , -0.975            // 1978
        , -1.152    , -0.975            // 1979
        , -0.797    , -0.797            // 1980
        , -0.975    , -0.797            // 1981
        , -0.797    , -0.975            // 1982
        , -0.975    , -0.975            // 1983
        , -2.747    , -0.089            // 1984
        , -2.569    , -0.089            // 1985
        , -2.747    , -0.266            // 1986
        , -2.569    , -0.266            // 1987
        , -2.215    , -0.089            // 1988
        , -2.392    , -0.089            // 1989
        , -2.215    , -0.266            // 1990
        , -2.392    , -0.266            // 1991
        , -2.747    ,  -0.62            // 1992
        , -2.569    ,  -0.62            // 1993
        , -2.747    , -0.443            // 1994
        , -2.569    , -0.443            // 1995
        , -2.215    ,  -0.62            // 1996
        , -2.392    ,  -0.62            // 1997
        , -2.215    , -0.443            // 1998
        , -2.392    , -0.443            // 1999
        , -1.506    , -0.089            // 2000
        , -1.683    , -0.089            // 2001
        , -1.506    , -0.266            // 2002
        , -1.683    , -0.266            // 2003
        , -2.038    , -0.089            // 2004
        , -1.861    , -0.089            // 2005
        , -2.038    , -0.266            // 2006
        , -1.861    , -0.266            // 2007
        , -1.506    ,  -0.62            // 2008
        , -1.683    ,  -0.62            // 2009
        , -1.506    , -0.443            // 2010
        , -1.683    , -0.443            // 2011
        , -2.038    ,  -0.62            // 2012
        , -1.861    ,  -0.62            // 2013
        , -2.038    , -0.443            // 2014
        , -1.861    , -0.443            // 2015
        , -2.747    , -1.329            // 2016
        , -2.569    , -1.329            // 2017
        , -2.747    , -1.152            // 2018
        , -2.569    , -1.152            // 2019
        , -2.215    , -1.329            // 2020
        , -2.392    , -1.329            // 2021
        , -2.215    , -1.152            // 2022
        , -2.392    , -1.152            // 2023
        , -2.747    , -0.797            // 2024
        , -2.569    , -0.797            // 2025
        , -2.747    , -0.975            // 2026
        , -2.569    , -0.975            // 2027
        , -2.215    , -0.797            // 2028
        , -2.392    , -0.797            // 2029
        , -2.215    , -0.975            // 2030
        , -2.392    , -0.975            // 2031
        , -1.506    , -1.329            // 2032
        , -1.683    , -1.329            // 2033
        , -1.506    , -1.152            // 2034
        , -1.683    , -1.152            // 2035
        , -2.038    , -1.329            // 2036
        , -1.861    , -1.329            // 2037
        , -2.038    , -1.152            // 2038
        , -1.861    , -1.152            // 2039
        , -1.506    , -0.797            // 2040
        , -1.683    , -0.797            // 2041
        , -1.506    , -0.975            // 2042
        , -1.683    , -0.975            // 2043
        , -2.038    , -0.797            // 2044
        , -1.861    , -0.797            // 2045
        , -2.038    , -0.975            // 2046
        , -1.861    , -0.975            // 2047
    };