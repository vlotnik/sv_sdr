    DVBS2X_APSK8_L_26_45 : super.plane = {
          -0.165    ,      0            // 0
        , -0.473    , -0.943            // 1
        , -0.473    ,  0.943            // 2
        , -1.322    ,      0            // 3
        ,  0.165    ,      0            // 4
        ,  0.473    , -0.943            // 5
        ,  0.473    ,  0.943            // 6
        ,  1.322    ,      0            // 7
    };