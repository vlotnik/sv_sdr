    //      I           Q
    GFSK2 : super.plane = {
           1.000    ,  0.000            // 0
        , -1.000    ,  0.000            // 1
    };