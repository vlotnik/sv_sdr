//--------------------------------------------------------------------------------------------------------------------------------
// name : raxi_bfm
//--------------------------------------------------------------------------------------------------------------------------------
interface raxi_bfm #(
      DW = 8
    , UW = 8
    , IW = 8
) (
      input                             clk
);
//--------------------------------------------------------------------------------------------------------------------------------
    bit                                 reset;
    bit                                 valid;
    bit                                 first;
    bit                                 last;
    bit                                 keep;
    bit                                 ready;
    bit[DW-1:0]                         data;
    bit[UW-1:0]                         user;
    bit[IW-1:0]                         id;

//--------------------------------------------------------------------------------------------------------------------------------
endinterface