    DVBS2_APSK16_4_5 : super.plane = {
           0.799    ,  0.799            // 0
        ,  0.799    , -0.799            // 1
        , -0.799    ,  0.799            // 2
        , -0.799    , -0.799            // 3
        ,  1.092    ,  0.292            // 4
        ,  1.092    , -0.292            // 5
        , -1.092    ,  0.292            // 6
        , -1.092    , -0.292            // 7
        ,  0.292    ,  1.092            // 8
        ,  0.292    , -1.092            // 9
        , -0.292    ,  1.092            // 10
        , -0.292    , -1.092            // 11
        ,  0.291    ,  0.291            // 12
        ,  0.291    , -0.291            // 13
        , -0.291    ,  0.291            // 14
        , -0.291    , -0.291            // 15
    };