    DVBS2_APSK32_4_5 : super.plane = {
           0.501    ,  0.501            // 0
        ,  0.183    ,  0.684            // 1
        ,  0.501    , -0.501            // 2
        ,  0.183    , -0.684            // 3
        , -0.501    ,  0.501            // 4
        , -0.183    ,  0.684            // 5
        , -0.501    , -0.501            // 6
        , -0.183    , -0.684            // 7
        ,  1.171    ,  0.485            // 8
        ,  0.485    ,  1.171            // 9
        ,  0.896    , -0.896            // 10
        ,      0    , -1.268            // 11
        , -0.896    ,  0.896            // 12
        ,      0    ,  1.268            // 13
        , -1.171    , -0.485            // 14
        , -0.485    , -1.171            // 15
        ,  0.684    ,  0.183            // 16
        ,  0.184    ,  0.184            // 17
        ,  0.684    , -0.183            // 18
        ,  0.184    , -0.184            // 19
        , -0.684    ,  0.183            // 20
        , -0.184    ,  0.184            // 21
        , -0.684    , -0.183            // 22
        , -0.184    , -0.184            // 23
        ,  1.268    ,      0            // 24
        ,  0.896    ,  0.896            // 25
        ,  1.171    , -0.485            // 26
        ,  0.485    , -1.171            // 27
        , -1.171    ,  0.485            // 28
        , -0.485    ,  1.171            // 29
        , -1.268    ,      0            // 30
        , -0.896    , -0.896            // 31
    };