    DVBS2_APSK16_5_6 : super.plane = {
           0.798    ,  0.798            // 0
        ,  0.798    , -0.798            // 1
        , -0.798    ,  0.798            // 2
        , -0.798    , -0.798            // 3
        ,  1.091    ,  0.292            // 4
        ,  1.091    , -0.292            // 5
        , -1.091    ,  0.292            // 6
        , -1.091    , -0.292            // 7
        ,  0.292    ,  1.091            // 8
        ,  0.292    , -1.091            // 9
        , -0.292    ,  1.091            // 10
        , -0.292    , -1.091            // 11
        ,  0.296    ,  0.296            // 12
        ,  0.296    , -0.296            // 13
        , -0.296    ,  0.296            // 14
        , -0.296    , -0.296            // 15
    };