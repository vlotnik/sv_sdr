    DVBS2X_4_12_16RBAPSK_2_3 : super.plane = {
          -0.715    ,  1.071            // 0
        , -0.251    ,  1.263            // 1
        ,  0.715    ,  1.071            // 2
        ,  0.251    ,  1.263            // 3
        , -0.468    ,  0.468            // 4
        , -0.171    ,  0.639            // 5
        ,  0.468    ,  0.468            // 6
        ,  0.171    ,  0.639            // 7
        , -1.071    ,  0.715            // 8
        , -1.263    ,  0.251            // 9
        ,  1.071    ,  0.715            // 10
        ,  1.263    ,  0.251            // 11
        , -0.639    ,  0.171            // 12
        , -0.164    ,  0.164            // 13
        ,  0.639    ,  0.171            // 14
        ,  0.164    ,  0.164            // 15
        , -0.715    , -1.071            // 16
        , -0.251    , -1.263            // 17
        ,  0.715    , -1.071            // 18
        ,  0.251    , -1.263            // 19
        , -0.468    , -0.468            // 20
        , -0.171    , -0.639            // 21
        ,  0.468    , -0.468            // 22
        ,  0.171    , -0.639            // 23
        , -1.071    , -0.715            // 24
        , -1.263    , -0.251            // 25
        ,  1.071    , -0.715            // 26
        ,  1.263    , -0.251            // 27
        , -0.639    , -0.171            // 28
        , -0.164    , -0.164            // 29
        ,  0.639    , -0.171            // 30
        ,  0.164    , -0.164            // 31
    };