    QAM64 : super.plane = {
           1.231    ,  1.231            // 0
        ,  1.231    ,   0.88            // 1
        ,   0.88    ,  1.231            // 2
        ,   0.88    ,   0.88            // 3
        ,  1.231    ,  0.528            // 4
        ,  1.231    ,  0.176            // 5
        ,   0.88    ,  0.528            // 6
        ,   0.88    ,  0.176            // 7
        ,  0.528    ,  1.231            // 8
        ,  0.528    ,   0.88            // 9
        ,  0.176    ,  1.231            // 10
        ,  0.176    ,   0.88            // 11
        ,  0.528    ,  0.528            // 12
        ,  0.528    ,  0.176            // 13
        ,  0.176    ,  0.528            // 14
        ,  0.176    ,  0.176            // 15
        ,  1.231    , -0.176            // 16
        ,  1.231    , -0.528            // 17
        ,   0.88    , -0.176            // 18
        ,   0.88    , -0.528            // 19
        ,  1.231    ,  -0.88            // 20
        ,  1.231    , -1.231            // 21
        ,   0.88    ,  -0.88            // 22
        ,   0.88    , -1.231            // 23
        ,  0.528    , -0.176            // 24
        ,  0.528    , -0.528            // 25
        ,  0.176    , -0.176            // 26
        ,  0.176    , -0.528            // 27
        ,  0.528    ,  -0.88            // 28
        ,  0.528    , -1.231            // 29
        ,  0.176    ,  -0.88            // 30
        ,  0.176    , -1.231            // 31
        , -0.176    ,  1.231            // 32
        , -0.176    ,   0.88            // 33
        , -0.528    ,  1.231            // 34
        , -0.528    ,   0.88            // 35
        , -0.176    ,  0.528            // 36
        , -0.176    ,  0.176            // 37
        , -0.528    ,  0.528            // 38
        , -0.528    ,  0.176            // 39
        ,  -0.88    ,  1.231            // 40
        ,  -0.88    ,   0.88            // 41
        , -1.231    ,  1.231            // 42
        , -1.231    ,   0.88            // 43
        ,  -0.88    ,  0.528            // 44
        ,  -0.88    ,  0.176            // 45
        , -1.231    ,  0.528            // 46
        , -1.231    ,  0.176            // 47
        , -0.176    , -0.176            // 48
        , -0.176    , -0.528            // 49
        , -0.528    , -0.176            // 50
        , -0.528    , -0.528            // 51
        , -0.176    ,  -0.88            // 52
        , -0.176    , -1.231            // 53
        , -0.528    ,  -0.88            // 54
        , -0.528    , -1.231            // 55
        ,  -0.88    , -0.176            // 56
        ,  -0.88    , -0.528            // 57
        , -1.231    , -0.176            // 58
        , -1.231    , -0.528            // 59
        ,  -0.88    ,  -0.88            // 60
        ,  -0.88    , -1.231            // 61
        , -1.231    ,  -0.88            // 62
        , -1.231    , -1.231            // 63
    };