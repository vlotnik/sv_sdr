    DVBS2_APSK32_3_4 : super.plane = {
           0.487    ,  0.487            // 0
        ,  0.178    ,  0.665            // 1
        ,  0.487    , -0.487            // 2
        ,  0.178    , -0.665            // 3
        , -0.487    ,  0.487            // 4
        , -0.178    ,  0.665            // 5
        , -0.487    , -0.487            // 6
        , -0.178    , -0.665            // 7
        ,   1.18    ,  0.489            // 8
        ,  0.489    ,   1.18            // 9
        ,  0.903    , -0.903            // 10
        ,      0    , -1.277            // 11
        , -0.903    ,  0.903            // 12
        ,      0    ,  1.277            // 13
        ,  -1.18    , -0.489            // 14
        , -0.489    ,  -1.18            // 15
        ,  0.665    ,  0.178            // 16
        ,  0.171    ,  0.171            // 17
        ,  0.665    , -0.178            // 18
        ,  0.171    , -0.171            // 19
        , -0.665    ,  0.178            // 20
        , -0.171    ,  0.171            // 21
        , -0.665    , -0.178            // 22
        , -0.171    , -0.171            // 23
        ,  1.277    ,      0            // 24
        ,  0.903    ,  0.903            // 25
        ,   1.18    , -0.489            // 26
        ,  0.489    ,  -1.18            // 27
        ,  -1.18    ,  0.489            // 28
        , -0.489    ,   1.18            // 29
        , -1.277    ,      0            // 30
        , -0.903    , -0.903            // 31
    };