    DVBS2_APSK32_9_10 : super.plane = {
           0.521    ,  0.521            // 0
        ,  0.191    ,  0.712            // 1
        ,  0.521    , -0.521            // 2
        ,  0.191    , -0.712            // 3
        , -0.521    ,  0.521            // 4
        , -0.191    ,  0.712            // 5
        , -0.521    , -0.521            // 6
        , -0.191    , -0.712            // 7
        ,  1.158    ,   0.48            // 8
        ,   0.48    ,  1.158            // 9
        ,  0.886    , -0.886            // 10
        ,      0    , -1.253            // 11
        , -0.886    ,  0.886            // 12
        ,      0    ,  1.253            // 13
        , -1.158    ,  -0.48            // 14
        ,  -0.48    , -1.158            // 15
        ,  0.712    ,  0.191            // 16
        ,  0.206    ,  0.206            // 17
        ,  0.712    , -0.191            // 18
        ,  0.206    , -0.206            // 19
        , -0.712    ,  0.191            // 20
        , -0.206    ,  0.206            // 21
        , -0.712    , -0.191            // 22
        , -0.206    , -0.206            // 23
        ,  1.253    ,      0            // 24
        ,  0.886    ,  0.886            // 25
        ,  1.158    ,  -0.48            // 26
        ,   0.48    , -1.158            // 27
        , -1.158    ,   0.48            // 28
        ,  -0.48    ,  1.158            // 29
        , -1.253    ,      0            // 30
        , -0.886    , -0.886            // 31
    };