    DVBS2X_4_8_4_16APSK_128_180 : super.plane = {
           0.164    ,  0.164            // 0
        ,  0.253    ,  1.274            // 1
        ,  0.164    , -0.164            // 2
        ,  0.253    , -1.274            // 3
        , -0.164    ,  0.164            // 4
        , -0.253    ,  1.274            // 5
        , -0.164    , -0.164            // 6
        , -0.253    , -1.274            // 7
        ,  0.582    ,  0.156            // 8
        ,  1.274    ,  0.253            // 9
        ,  0.582    , -0.156            // 10
        ,  1.274    , -0.253            // 11
        , -0.582    ,  0.156            // 12
        , -1.274    ,  0.253            // 13
        , -0.582    , -0.156            // 14
        , -1.274    , -0.253            // 15
        ,  0.156    ,  0.582            // 16
        ,  0.721    ,   1.08            // 17
        ,  0.156    , -0.582            // 18
        ,  0.721    ,  -1.08            // 19
        , -0.156    ,  0.582            // 20
        , -0.721    ,   1.08            // 21
        , -0.156    , -0.582            // 22
        , -0.721    ,  -1.08            // 23
        ,   0.49    ,   0.49            // 24
        ,   1.08    ,  0.721            // 25
        ,   0.49    ,  -0.49            // 26
        ,   1.08    , -0.721            // 27
        ,  -0.49    ,   0.49            // 28
        ,  -1.08    ,  0.721            // 29
        ,  -0.49    ,  -0.49            // 30
        ,  -1.08    , -0.721            // 31
    };