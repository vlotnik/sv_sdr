    QAM16, QAM16_POL : super.plane = {
           1.061    ,  1.061            // 0
        ,  1.061    ,  0.354            // 1
        ,  0.354    ,  1.061            // 2
        ,  0.354    ,  0.354            // 3
        ,  1.061    , -0.354            // 4
        ,  1.061    , -1.061            // 5
        ,  0.354    , -0.354            // 6
        ,  0.354    , -1.061            // 7
        , -0.354    ,  1.061            // 8
        , -0.354    ,  0.354            // 9
        , -1.061    ,  1.061            // 10
        , -1.061    ,  0.354            // 11
        , -0.354    , -0.354            // 12
        , -0.354    , -1.061            // 13
        , -1.061    , -0.354            // 14
        , -1.061    , -1.061            // 15
    };