    DVBS2X_256APSK_135_180 : super.plane = {
           0.288    ,  0.028            // 0
        ,  0.277    ,  0.084            // 1
        ,  0.224    ,  0.184            // 2
        ,  0.255    ,  0.137            // 3
        ,  0.028    ,  0.288            // 4
        ,  0.084    ,  0.277            // 5
        ,  0.184    ,  0.224            // 6
        ,  0.137    ,  0.255            // 7
        , -0.288    ,  0.028            // 8
        , -0.277    ,  0.084            // 9
        , -0.224    ,  0.184            // 10
        , -0.255    ,  0.137            // 11
        , -0.028    ,  0.288            // 12
        , -0.084    ,  0.277            // 13
        , -0.184    ,  0.224            // 14
        , -0.137    ,  0.255            // 15
        ,  0.288    , -0.028            // 16
        ,  0.277    , -0.084            // 17
        ,  0.224    , -0.184            // 18
        ,  0.255    , -0.137            // 19
        ,  0.028    , -0.288            // 20
        ,  0.084    , -0.277            // 21
        ,  0.184    , -0.224            // 22
        ,  0.137    , -0.255            // 23
        , -0.288    , -0.028            // 24
        , -0.277    , -0.084            // 25
        , -0.224    , -0.184            // 26
        , -0.255    , -0.137            // 27
        , -0.028    , -0.288            // 28
        , -0.084    , -0.277            // 29
        , -0.184    , -0.224            // 30
        , -0.137    , -0.255            // 31
        ,  0.517    ,  0.051            // 32
        ,  0.497    ,  0.151            // 33
        ,  0.402    ,   0.33            // 34
        ,  0.458    ,  0.245            // 35
        ,  0.051    ,  0.517            // 36
        ,  0.151    ,  0.497            // 37
        ,   0.33    ,  0.402            // 38
        ,  0.245    ,  0.458            // 39
        , -0.517    ,  0.051            // 40
        , -0.497    ,  0.151            // 41
        , -0.402    ,   0.33            // 42
        , -0.458    ,  0.245            // 43
        , -0.051    ,  0.517            // 44
        , -0.151    ,  0.497            // 45
        ,  -0.33    ,  0.402            // 46
        , -0.245    ,  0.458            // 47
        ,  0.517    , -0.051            // 48
        ,  0.497    , -0.151            // 49
        ,  0.402    ,  -0.33            // 50
        ,  0.458    , -0.245            // 51
        ,  0.051    , -0.517            // 52
        ,  0.151    , -0.497            // 53
        ,   0.33    , -0.402            // 54
        ,  0.245    , -0.458            // 55
        , -0.517    , -0.051            // 56
        , -0.497    , -0.151            // 57
        , -0.402    ,  -0.33            // 58
        , -0.458    , -0.245            // 59
        , -0.051    , -0.517            // 60
        , -0.151    , -0.497            // 61
        ,  -0.33    , -0.402            // 62
        , -0.245    , -0.458            // 63
        ,  0.861    ,  0.085            // 64
        ,  0.828    ,  0.251            // 65
        ,  0.668    ,  0.549            // 66
        ,  0.763    ,  0.408            // 67
        ,  0.085    ,  0.861            // 68
        ,  0.251    ,  0.828            // 69
        ,  0.549    ,  0.668            // 70
        ,  0.408    ,  0.763            // 71
        , -0.861    ,  0.085            // 72
        , -0.828    ,  0.251            // 73
        , -0.668    ,  0.549            // 74
        , -0.763    ,  0.408            // 75
        , -0.085    ,  0.861            // 76
        , -0.251    ,  0.828            // 77
        , -0.549    ,  0.668            // 78
        , -0.408    ,  0.763            // 79
        ,  0.861    , -0.085            // 80
        ,  0.828    , -0.251            // 81
        ,  0.668    , -0.549            // 82
        ,  0.763    , -0.408            // 83
        ,  0.085    , -0.861            // 84
        ,  0.251    , -0.828            // 85
        ,  0.549    , -0.668            // 86
        ,  0.408    , -0.763            // 87
        , -0.861    , -0.085            // 88
        , -0.828    , -0.251            // 89
        , -0.668    , -0.549            // 90
        , -0.763    , -0.408            // 91
        , -0.085    , -0.861            // 92
        , -0.251    , -0.828            // 93
        , -0.549    , -0.668            // 94
        , -0.408    , -0.763            // 95
        ,  0.694    ,  0.068            // 96
        ,  0.668    ,  0.203            // 97
        ,  0.539    ,  0.443            // 98
        ,  0.615    ,  0.329            // 99
        ,  0.068    ,  0.694            // 100
        ,  0.203    ,  0.668            // 101
        ,  0.443    ,  0.539            // 102
        ,  0.329    ,  0.615            // 103
        , -0.694    ,  0.068            // 104
        , -0.668    ,  0.203            // 105
        , -0.539    ,  0.443            // 106
        , -0.615    ,  0.329            // 107
        , -0.068    ,  0.694            // 108
        , -0.203    ,  0.668            // 109
        , -0.443    ,  0.539            // 110
        , -0.329    ,  0.615            // 111
        ,  0.694    , -0.068            // 112
        ,  0.668    , -0.203            // 113
        ,  0.539    , -0.443            // 114
        ,  0.615    , -0.329            // 115
        ,  0.068    , -0.694            // 116
        ,  0.203    , -0.668            // 117
        ,  0.443    , -0.539            // 118
        ,  0.329    , -0.615            // 119
        , -0.694    , -0.068            // 120
        , -0.668    , -0.203            // 121
        , -0.539    , -0.443            // 122
        , -0.615    , -0.329            // 123
        , -0.068    , -0.694            // 124
        , -0.203    , -0.668            // 125
        , -0.443    , -0.539            // 126
        , -0.329    , -0.615            // 127
        ,  1.499    ,  0.148            // 128
        ,  1.441    ,  0.437            // 129
        ,  1.164    ,  0.955            // 130
        ,  1.328    ,   0.71            // 131
        ,  0.148    ,  1.499            // 132
        ,  0.437    ,  1.441            // 133
        ,  0.955    ,  1.164            // 134
        ,   0.71    ,  1.328            // 135
        , -1.499    ,  0.148            // 136
        , -1.441    ,  0.437            // 137
        , -1.164    ,  0.955            // 138
        , -1.328    ,   0.71            // 139
        , -0.148    ,  1.499            // 140
        , -0.437    ,  1.441            // 141
        , -0.955    ,  1.164            // 142
        ,  -0.71    ,  1.328            // 143
        ,  1.499    , -0.148            // 144
        ,  1.441    , -0.437            // 145
        ,  1.164    , -0.955            // 146
        ,  1.328    ,  -0.71            // 147
        ,  0.148    , -1.499            // 148
        ,  0.437    , -1.441            // 149
        ,  0.955    , -1.164            // 150
        ,   0.71    , -1.328            // 151
        , -1.499    , -0.148            // 152
        , -1.441    , -0.437            // 153
        , -1.164    , -0.955            // 154
        , -1.328    ,  -0.71            // 155
        , -0.148    , -1.499            // 156
        , -0.437    , -1.441            // 157
        , -0.955    , -1.164            // 158
        ,  -0.71    , -1.328            // 159
        ,  1.297    ,  0.128            // 160
        ,  1.247    ,  0.378            // 161
        ,  1.007    ,  0.827            // 162
        ,  1.149    ,  0.614            // 163
        ,  0.128    ,  1.297            // 164
        ,  0.378    ,  1.247            // 165
        ,  0.827    ,  1.007            // 166
        ,  0.614    ,  1.149            // 167
        , -1.297    ,  0.128            // 168
        , -1.247    ,  0.378            // 169
        , -1.007    ,  0.827            // 170
        , -1.149    ,  0.614            // 171
        , -0.128    ,  1.297            // 172
        , -0.378    ,  1.247            // 173
        , -0.827    ,  1.007            // 174
        , -0.614    ,  1.149            // 175
        ,  1.297    , -0.128            // 176
        ,  1.247    , -0.378            // 177
        ,  1.007    , -0.827            // 178
        ,  1.149    , -0.614            // 179
        ,  0.128    , -1.297            // 180
        ,  0.378    , -1.247            // 181
        ,  0.827    , -1.007            // 182
        ,  0.614    , -1.149            // 183
        , -1.297    , -0.128            // 184
        , -1.247    , -0.378            // 185
        , -1.007    , -0.827            // 186
        , -1.149    , -0.614            // 187
        , -0.128    , -1.297            // 188
        , -0.378    , -1.247            // 189
        , -0.827    , -1.007            // 190
        , -0.614    , -1.149            // 191
        ,  1.031    ,  0.102            // 192
        ,  0.992    ,  0.301            // 193
        ,  0.801    ,  0.658            // 194
        ,  0.914    ,  0.489            // 195
        ,  0.102    ,  1.031            // 196
        ,  0.301    ,  0.992            // 197
        ,  0.658    ,  0.801            // 198
        ,  0.489    ,  0.914            // 199
        , -1.031    ,  0.102            // 200
        , -0.992    ,  0.301            // 201
        , -0.801    ,  0.658            // 202
        , -0.914    ,  0.489            // 203
        , -0.102    ,  1.031            // 204
        , -0.301    ,  0.992            // 205
        , -0.658    ,  0.801            // 206
        , -0.489    ,  0.914            // 207
        ,  1.031    , -0.102            // 208
        ,  0.992    , -0.301            // 209
        ,  0.801    , -0.658            // 210
        ,  0.914    , -0.489            // 211
        ,  0.102    , -1.031            // 212
        ,  0.301    , -0.992            // 213
        ,  0.658    , -0.801            // 214
        ,  0.489    , -0.914            // 215
        , -1.031    , -0.102            // 216
        , -0.992    , -0.301            // 217
        , -0.801    , -0.658            // 218
        , -0.914    , -0.489            // 219
        , -0.102    , -1.031            // 220
        , -0.301    , -0.992            // 221
        , -0.658    , -0.801            // 222
        , -0.489    , -0.914            // 223
        ,  1.166    ,  0.115            // 224
        ,  1.121    ,   0.34            // 225
        ,  0.906    ,  0.743            // 226
        ,  1.033    ,  0.552            // 227
        ,  0.115    ,  1.166            // 228
        ,   0.34    ,  1.121            // 229
        ,  0.743    ,  0.906            // 230
        ,  0.552    ,  1.033            // 231
        , -1.166    ,  0.115            // 232
        , -1.121    ,   0.34            // 233
        , -0.906    ,  0.743            // 234
        , -1.033    ,  0.552            // 235
        , -0.115    ,  1.166            // 236
        ,  -0.34    ,  1.121            // 237
        , -0.743    ,  0.906            // 238
        , -0.552    ,  1.033            // 239
        ,  1.166    , -0.115            // 240
        ,  1.121    ,  -0.34            // 241
        ,  0.906    , -0.743            // 242
        ,  1.033    , -0.552            // 243
        ,  0.115    , -1.166            // 244
        ,   0.34    , -1.121            // 245
        ,  0.743    , -0.906            // 246
        ,  0.552    , -1.033            // 247
        , -1.166    , -0.115            // 248
        , -1.121    ,  -0.34            // 249
        , -0.906    , -0.743            // 250
        , -1.033    , -0.552            // 251
        , -0.115    , -1.166            // 252
        ,  -0.34    , -1.121            // 253
        , -0.743    , -0.906            // 254
        , -0.552    , -1.033            // 255
    };