    DVBS2X_16_16_16_16APSK_128_180 : super.plane = {
           0.374    ,  0.074            // 0
        ,  0.317    ,  0.212            // 1
        ,  0.074    ,  0.374            // 2
        ,  0.212    ,  0.317            // 3
        , -0.374    ,  0.074            // 4
        , -0.317    ,  0.212            // 5
        , -0.074    ,  0.374            // 6
        , -0.212    ,  0.317            // 7
        ,  0.374    , -0.074            // 8
        ,  0.317    , -0.212            // 9
        ,  0.074    , -0.374            // 10
        ,  0.212    , -0.317            // 11
        , -0.374    , -0.074            // 12
        , -0.317    , -0.212            // 13
        , -0.074    , -0.374            // 14
        , -0.212    , -0.317            // 15
        ,  0.703    ,   0.14            // 16
        ,  0.596    ,  0.398            // 17
        ,   0.14    ,  0.703            // 18
        ,  0.398    ,  0.596            // 19
        , -0.703    ,   0.14            // 20
        , -0.596    ,  0.398            // 21
        ,  -0.14    ,  0.703            // 22
        , -0.398    ,  0.596            // 23
        ,  0.703    ,  -0.14            // 24
        ,  0.596    , -0.398            // 25
        ,   0.14    , -0.703            // 26
        ,  0.398    , -0.596            // 27
        , -0.703    ,  -0.14            // 28
        , -0.596    , -0.398            // 29
        ,  -0.14    , -0.703            // 30
        , -0.398    , -0.596            // 31
        ,  1.476    ,  0.294            // 32
        ,  1.252    ,  0.836            // 33
        ,  0.294    ,  1.476            // 34
        ,  0.836    ,  1.252            // 35
        , -1.476    ,  0.294            // 36
        , -1.252    ,  0.836            // 37
        , -0.294    ,  1.476            // 38
        , -0.836    ,  1.252            // 39
        ,  1.476    , -0.294            // 40
        ,  1.252    , -0.836            // 41
        ,  0.294    , -1.476            // 42
        ,  0.836    , -1.252            // 43
        , -1.476    , -0.294            // 44
        , -1.252    , -0.836            // 45
        , -0.294    , -1.476            // 46
        , -0.836    , -1.252            // 47
        ,  1.017    ,  0.202            // 48
        ,  0.862    ,  0.576            // 49
        ,  0.202    ,  1.017            // 50
        ,  0.576    ,  0.862            // 51
        , -1.017    ,  0.202            // 52
        , -0.862    ,  0.576            // 53
        , -0.202    ,  1.017            // 54
        , -0.576    ,  0.862            // 55
        ,  1.017    , -0.202            // 56
        ,  0.862    , -0.576            // 57
        ,  0.202    , -1.017            // 58
        ,  0.576    , -0.862            // 59
        , -1.017    , -0.202            // 60
        , -0.862    , -0.576            // 61
        , -0.202    , -1.017            // 62
        , -0.576    , -0.862            // 63
    };