    DVBS2X_4_12APSK_140_180 : super.plane = {
           0.806    ,  0.806            // 0
        ,  0.806    , -0.806            // 1
        , -0.806    ,  0.806            // 2
        , -0.806    , -0.806            // 3
        ,  1.101    ,  0.295            // 4
        ,  1.101    , -0.295            // 5
        , -1.101    ,  0.295            // 6
        , -1.101    , -0.295            // 7
        ,  0.295    ,  1.101            // 8
        ,  0.295    , -1.101            // 9
        , -0.295    ,  1.101            // 10
        , -0.295    , -1.101            // 11
        ,  0.224    ,  0.224            // 12
        ,  0.224    , -0.224            // 13
        , -0.224    ,  0.224            // 14
        , -0.224    , -0.224            // 15
    };