    QAM1024 : super.plane = {
           2.747    ,  2.747            // 0
        ,  2.747    ,  2.569            // 1
        ,  2.569    ,  2.747            // 2
        ,  2.569    ,  2.569            // 3
        ,  2.747    ,  2.392            // 4
        ,  2.747    ,  2.215            // 5
        ,  2.569    ,  2.392            // 6
        ,  2.569    ,  2.215            // 7
        ,  2.392    ,  2.747            // 8
        ,  2.392    ,  2.569            // 9
        ,  2.215    ,  2.747            // 10
        ,  2.215    ,  2.569            // 11
        ,  2.392    ,  2.392            // 12
        ,  2.392    ,  2.215            // 13
        ,  2.215    ,  2.392            // 14
        ,  2.215    ,  2.215            // 15
        ,  2.747    ,  2.038            // 16
        ,  2.747    ,  1.861            // 17
        ,  2.569    ,  2.038            // 18
        ,  2.569    ,  1.861            // 19
        ,  2.747    ,  1.683            // 20
        ,  2.747    ,  1.506            // 21
        ,  2.569    ,  1.683            // 22
        ,  2.569    ,  1.506            // 23
        ,  2.392    ,  2.038            // 24
        ,  2.392    ,  1.861            // 25
        ,  2.215    ,  2.038            // 26
        ,  2.215    ,  1.861            // 27
        ,  2.392    ,  1.683            // 28
        ,  2.392    ,  1.506            // 29
        ,  2.215    ,  1.683            // 30
        ,  2.215    ,  1.506            // 31
        ,  2.038    ,  2.747            // 32
        ,  2.038    ,  2.569            // 33
        ,  1.861    ,  2.747            // 34
        ,  1.861    ,  2.569            // 35
        ,  2.038    ,  2.392            // 36
        ,  2.038    ,  2.215            // 37
        ,  1.861    ,  2.392            // 38
        ,  1.861    ,  2.215            // 39
        ,  1.683    ,  2.747            // 40
        ,  1.683    ,  2.569            // 41
        ,  1.506    ,  2.747            // 42
        ,  1.506    ,  2.569            // 43
        ,  1.683    ,  2.392            // 44
        ,  1.683    ,  2.215            // 45
        ,  1.506    ,  2.392            // 46
        ,  1.506    ,  2.215            // 47
        ,  2.038    ,  2.038            // 48
        ,  2.038    ,  1.861            // 49
        ,  1.861    ,  2.038            // 50
        ,  1.861    ,  1.861            // 51
        ,  2.038    ,  1.683            // 52
        ,  2.038    ,  1.506            // 53
        ,  1.861    ,  1.683            // 54
        ,  1.861    ,  1.506            // 55
        ,  1.683    ,  2.038            // 56
        ,  1.683    ,  1.861            // 57
        ,  1.506    ,  2.038            // 58
        ,  1.506    ,  1.861            // 59
        ,  1.683    ,  1.683            // 60
        ,  1.683    ,  1.506            // 61
        ,  1.506    ,  1.683            // 62
        ,  1.506    ,  1.506            // 63
        ,  2.747    ,  1.329            // 64
        ,  2.747    ,  1.152            // 65
        ,  2.569    ,  1.329            // 66
        ,  2.569    ,  1.152            // 67
        ,  2.747    ,  0.975            // 68
        ,  2.747    ,  0.797            // 69
        ,  2.569    ,  0.975            // 70
        ,  2.569    ,  0.797            // 71
        ,  2.392    ,  1.329            // 72
        ,  2.392    ,  1.152            // 73
        ,  2.215    ,  1.329            // 74
        ,  2.215    ,  1.152            // 75
        ,  2.392    ,  0.975            // 76
        ,  2.392    ,  0.797            // 77
        ,  2.215    ,  0.975            // 78
        ,  2.215    ,  0.797            // 79
        ,  2.747    ,   0.62            // 80
        ,  2.747    ,  0.443            // 81
        ,  2.569    ,   0.62            // 82
        ,  2.569    ,  0.443            // 83
        ,  2.747    ,  0.266            // 84
        ,  2.747    ,  0.089            // 85
        ,  2.569    ,  0.266            // 86
        ,  2.569    ,  0.089            // 87
        ,  2.392    ,   0.62            // 88
        ,  2.392    ,  0.443            // 89
        ,  2.215    ,   0.62            // 90
        ,  2.215    ,  0.443            // 91
        ,  2.392    ,  0.266            // 92
        ,  2.392    ,  0.089            // 93
        ,  2.215    ,  0.266            // 94
        ,  2.215    ,  0.089            // 95
        ,  2.038    ,  1.329            // 96
        ,  2.038    ,  1.152            // 97
        ,  1.861    ,  1.329            // 98
        ,  1.861    ,  1.152            // 99
        ,  2.038    ,  0.975            // 100
        ,  2.038    ,  0.797            // 101
        ,  1.861    ,  0.975            // 102
        ,  1.861    ,  0.797            // 103
        ,  1.683    ,  1.329            // 104
        ,  1.683    ,  1.152            // 105
        ,  1.506    ,  1.329            // 106
        ,  1.506    ,  1.152            // 107
        ,  1.683    ,  0.975            // 108
        ,  1.683    ,  0.797            // 109
        ,  1.506    ,  0.975            // 110
        ,  1.506    ,  0.797            // 111
        ,  2.038    ,   0.62            // 112
        ,  2.038    ,  0.443            // 113
        ,  1.861    ,   0.62            // 114
        ,  1.861    ,  0.443            // 115
        ,  2.038    ,  0.266            // 116
        ,  2.038    ,  0.089            // 117
        ,  1.861    ,  0.266            // 118
        ,  1.861    ,  0.089            // 119
        ,  1.683    ,   0.62            // 120
        ,  1.683    ,  0.443            // 121
        ,  1.506    ,   0.62            // 122
        ,  1.506    ,  0.443            // 123
        ,  1.683    ,  0.266            // 124
        ,  1.683    ,  0.089            // 125
        ,  1.506    ,  0.266            // 126
        ,  1.506    ,  0.089            // 127
        ,  1.329    ,  2.747            // 128
        ,  1.329    ,  2.569            // 129
        ,  1.152    ,  2.747            // 130
        ,  1.152    ,  2.569            // 131
        ,  1.329    ,  2.392            // 132
        ,  1.329    ,  2.215            // 133
        ,  1.152    ,  2.392            // 134
        ,  1.152    ,  2.215            // 135
        ,  0.975    ,  2.747            // 136
        ,  0.975    ,  2.569            // 137
        ,  0.797    ,  2.747            // 138
        ,  0.797    ,  2.569            // 139
        ,  0.975    ,  2.392            // 140
        ,  0.975    ,  2.215            // 141
        ,  0.797    ,  2.392            // 142
        ,  0.797    ,  2.215            // 143
        ,  1.329    ,  2.038            // 144
        ,  1.329    ,  1.861            // 145
        ,  1.152    ,  2.038            // 146
        ,  1.152    ,  1.861            // 147
        ,  1.329    ,  1.683            // 148
        ,  1.329    ,  1.506            // 149
        ,  1.152    ,  1.683            // 150
        ,  1.152    ,  1.506            // 151
        ,  0.975    ,  2.038            // 152
        ,  0.975    ,  1.861            // 153
        ,  0.797    ,  2.038            // 154
        ,  0.797    ,  1.861            // 155
        ,  0.975    ,  1.683            // 156
        ,  0.975    ,  1.506            // 157
        ,  0.797    ,  1.683            // 158
        ,  0.797    ,  1.506            // 159
        ,   0.62    ,  2.747            // 160
        ,   0.62    ,  2.569            // 161
        ,  0.443    ,  2.747            // 162
        ,  0.443    ,  2.569            // 163
        ,   0.62    ,  2.392            // 164
        ,   0.62    ,  2.215            // 165
        ,  0.443    ,  2.392            // 166
        ,  0.443    ,  2.215            // 167
        ,  0.266    ,  2.747            // 168
        ,  0.266    ,  2.569            // 169
        ,  0.089    ,  2.747            // 170
        ,  0.089    ,  2.569            // 171
        ,  0.266    ,  2.392            // 172
        ,  0.266    ,  2.215            // 173
        ,  0.089    ,  2.392            // 174
        ,  0.089    ,  2.215            // 175
        ,   0.62    ,  2.038            // 176
        ,   0.62    ,  1.861            // 177
        ,  0.443    ,  2.038            // 178
        ,  0.443    ,  1.861            // 179
        ,   0.62    ,  1.683            // 180
        ,   0.62    ,  1.506            // 181
        ,  0.443    ,  1.683            // 182
        ,  0.443    ,  1.506            // 183
        ,  0.266    ,  2.038            // 184
        ,  0.266    ,  1.861            // 185
        ,  0.089    ,  2.038            // 186
        ,  0.089    ,  1.861            // 187
        ,  0.266    ,  1.683            // 188
        ,  0.266    ,  1.506            // 189
        ,  0.089    ,  1.683            // 190
        ,  0.089    ,  1.506            // 191
        ,  1.329    ,  1.329            // 192
        ,  1.329    ,  1.152            // 193
        ,  1.152    ,  1.329            // 194
        ,  1.152    ,  1.152            // 195
        ,  1.329    ,  0.975            // 196
        ,  1.329    ,  0.797            // 197
        ,  1.152    ,  0.975            // 198
        ,  1.152    ,  0.797            // 199
        ,  0.975    ,  1.329            // 200
        ,  0.975    ,  1.152            // 201
        ,  0.797    ,  1.329            // 202
        ,  0.797    ,  1.152            // 203
        ,  0.975    ,  0.975            // 204
        ,  0.975    ,  0.797            // 205
        ,  0.797    ,  0.975            // 206
        ,  0.797    ,  0.797            // 207
        ,  1.329    ,   0.62            // 208
        ,  1.329    ,  0.443            // 209
        ,  1.152    ,   0.62            // 210
        ,  1.152    ,  0.443            // 211
        ,  1.329    ,  0.266            // 212
        ,  1.329    ,  0.089            // 213
        ,  1.152    ,  0.266            // 214
        ,  1.152    ,  0.089            // 215
        ,  0.975    ,   0.62            // 216
        ,  0.975    ,  0.443            // 217
        ,  0.797    ,   0.62            // 218
        ,  0.797    ,  0.443            // 219
        ,  0.975    ,  0.266            // 220
        ,  0.975    ,  0.089            // 221
        ,  0.797    ,  0.266            // 222
        ,  0.797    ,  0.089            // 223
        ,   0.62    ,  1.329            // 224
        ,   0.62    ,  1.152            // 225
        ,  0.443    ,  1.329            // 226
        ,  0.443    ,  1.152            // 227
        ,   0.62    ,  0.975            // 228
        ,   0.62    ,  0.797            // 229
        ,  0.443    ,  0.975            // 230
        ,  0.443    ,  0.797            // 231
        ,  0.266    ,  1.329            // 232
        ,  0.266    ,  1.152            // 233
        ,  0.089    ,  1.329            // 234
        ,  0.089    ,  1.152            // 235
        ,  0.266    ,  0.975            // 236
        ,  0.266    ,  0.797            // 237
        ,  0.089    ,  0.975            // 238
        ,  0.089    ,  0.797            // 239
        ,   0.62    ,   0.62            // 240
        ,   0.62    ,  0.443            // 241
        ,  0.443    ,   0.62            // 242
        ,  0.443    ,  0.443            // 243
        ,   0.62    ,  0.266            // 244
        ,   0.62    ,  0.089            // 245
        ,  0.443    ,  0.266            // 246
        ,  0.443    ,  0.089            // 247
        ,  0.266    ,   0.62            // 248
        ,  0.266    ,  0.443            // 249
        ,  0.089    ,   0.62            // 250
        ,  0.089    ,  0.443            // 251
        ,  0.266    ,  0.266            // 252
        ,  0.266    ,  0.089            // 253
        ,  0.089    ,  0.266            // 254
        ,  0.089    ,  0.089            // 255
        ,  2.747    , -0.089            // 256
        ,  2.747    , -0.266            // 257
        ,  2.569    , -0.089            // 258
        ,  2.569    , -0.266            // 259
        ,  2.747    , -0.443            // 260
        ,  2.747    ,  -0.62            // 261
        ,  2.569    , -0.443            // 262
        ,  2.569    ,  -0.62            // 263
        ,  2.392    , -0.089            // 264
        ,  2.392    , -0.266            // 265
        ,  2.215    , -0.089            // 266
        ,  2.215    , -0.266            // 267
        ,  2.392    , -0.443            // 268
        ,  2.392    ,  -0.62            // 269
        ,  2.215    , -0.443            // 270
        ,  2.215    ,  -0.62            // 271
        ,  2.747    , -0.797            // 272
        ,  2.747    , -0.975            // 273
        ,  2.569    , -0.797            // 274
        ,  2.569    , -0.975            // 275
        ,  2.747    , -1.152            // 276
        ,  2.747    , -1.329            // 277
        ,  2.569    , -1.152            // 278
        ,  2.569    , -1.329            // 279
        ,  2.392    , -0.797            // 280
        ,  2.392    , -0.975            // 281
        ,  2.215    , -0.797            // 282
        ,  2.215    , -0.975            // 283
        ,  2.392    , -1.152            // 284
        ,  2.392    , -1.329            // 285
        ,  2.215    , -1.152            // 286
        ,  2.215    , -1.329            // 287
        ,  2.038    , -0.089            // 288
        ,  2.038    , -0.266            // 289
        ,  1.861    , -0.089            // 290
        ,  1.861    , -0.266            // 291
        ,  2.038    , -0.443            // 292
        ,  2.038    ,  -0.62            // 293
        ,  1.861    , -0.443            // 294
        ,  1.861    ,  -0.62            // 295
        ,  1.683    , -0.089            // 296
        ,  1.683    , -0.266            // 297
        ,  1.506    , -0.089            // 298
        ,  1.506    , -0.266            // 299
        ,  1.683    , -0.443            // 300
        ,  1.683    ,  -0.62            // 301
        ,  1.506    , -0.443            // 302
        ,  1.506    ,  -0.62            // 303
        ,  2.038    , -0.797            // 304
        ,  2.038    , -0.975            // 305
        ,  1.861    , -0.797            // 306
        ,  1.861    , -0.975            // 307
        ,  2.038    , -1.152            // 308
        ,  2.038    , -1.329            // 309
        ,  1.861    , -1.152            // 310
        ,  1.861    , -1.329            // 311
        ,  1.683    , -0.797            // 312
        ,  1.683    , -0.975            // 313
        ,  1.506    , -0.797            // 314
        ,  1.506    , -0.975            // 315
        ,  1.683    , -1.152            // 316
        ,  1.683    , -1.329            // 317
        ,  1.506    , -1.152            // 318
        ,  1.506    , -1.329            // 319
        ,  2.747    , -1.506            // 320
        ,  2.747    , -1.683            // 321
        ,  2.569    , -1.506            // 322
        ,  2.569    , -1.683            // 323
        ,  2.747    , -1.861            // 324
        ,  2.747    , -2.038            // 325
        ,  2.569    , -1.861            // 326
        ,  2.569    , -2.038            // 327
        ,  2.392    , -1.506            // 328
        ,  2.392    , -1.683            // 329
        ,  2.215    , -1.506            // 330
        ,  2.215    , -1.683            // 331
        ,  2.392    , -1.861            // 332
        ,  2.392    , -2.038            // 333
        ,  2.215    , -1.861            // 334
        ,  2.215    , -2.038            // 335
        ,  2.747    , -2.215            // 336
        ,  2.747    , -2.392            // 337
        ,  2.569    , -2.215            // 338
        ,  2.569    , -2.392            // 339
        ,  2.747    , -2.569            // 340
        ,  2.747    , -2.747            // 341
        ,  2.569    , -2.569            // 342
        ,  2.569    , -2.747            // 343
        ,  2.392    , -2.215            // 344
        ,  2.392    , -2.392            // 345
        ,  2.215    , -2.215            // 346
        ,  2.215    , -2.392            // 347
        ,  2.392    , -2.569            // 348
        ,  2.392    , -2.747            // 349
        ,  2.215    , -2.569            // 350
        ,  2.215    , -2.747            // 351
        ,  2.038    , -1.506            // 352
        ,  2.038    , -1.683            // 353
        ,  1.861    , -1.506            // 354
        ,  1.861    , -1.683            // 355
        ,  2.038    , -1.861            // 356
        ,  2.038    , -2.038            // 357
        ,  1.861    , -1.861            // 358
        ,  1.861    , -2.038            // 359
        ,  1.683    , -1.506            // 360
        ,  1.683    , -1.683            // 361
        ,  1.506    , -1.506            // 362
        ,  1.506    , -1.683            // 363
        ,  1.683    , -1.861            // 364
        ,  1.683    , -2.038            // 365
        ,  1.506    , -1.861            // 366
        ,  1.506    , -2.038            // 367
        ,  2.038    , -2.215            // 368
        ,  2.038    , -2.392            // 369
        ,  1.861    , -2.215            // 370
        ,  1.861    , -2.392            // 371
        ,  2.038    , -2.569            // 372
        ,  2.038    , -2.747            // 373
        ,  1.861    , -2.569            // 374
        ,  1.861    , -2.747            // 375
        ,  1.683    , -2.215            // 376
        ,  1.683    , -2.392            // 377
        ,  1.506    , -2.215            // 378
        ,  1.506    , -2.392            // 379
        ,  1.683    , -2.569            // 380
        ,  1.683    , -2.747            // 381
        ,  1.506    , -2.569            // 382
        ,  1.506    , -2.747            // 383
        ,  1.329    , -0.089            // 384
        ,  1.329    , -0.266            // 385
        ,  1.152    , -0.089            // 386
        ,  1.152    , -0.266            // 387
        ,  1.329    , -0.443            // 388
        ,  1.329    ,  -0.62            // 389
        ,  1.152    , -0.443            // 390
        ,  1.152    ,  -0.62            // 391
        ,  0.975    , -0.089            // 392
        ,  0.975    , -0.266            // 393
        ,  0.797    , -0.089            // 394
        ,  0.797    , -0.266            // 395
        ,  0.975    , -0.443            // 396
        ,  0.975    ,  -0.62            // 397
        ,  0.797    , -0.443            // 398
        ,  0.797    ,  -0.62            // 399
        ,  1.329    , -0.797            // 400
        ,  1.329    , -0.975            // 401
        ,  1.152    , -0.797            // 402
        ,  1.152    , -0.975            // 403
        ,  1.329    , -1.152            // 404
        ,  1.329    , -1.329            // 405
        ,  1.152    , -1.152            // 406
        ,  1.152    , -1.329            // 407
        ,  0.975    , -0.797            // 408
        ,  0.975    , -0.975            // 409
        ,  0.797    , -0.797            // 410
        ,  0.797    , -0.975            // 411
        ,  0.975    , -1.152            // 412
        ,  0.975    , -1.329            // 413
        ,  0.797    , -1.152            // 414
        ,  0.797    , -1.329            // 415
        ,   0.62    , -0.089            // 416
        ,   0.62    , -0.266            // 417
        ,  0.443    , -0.089            // 418
        ,  0.443    , -0.266            // 419
        ,   0.62    , -0.443            // 420
        ,   0.62    ,  -0.62            // 421
        ,  0.443    , -0.443            // 422
        ,  0.443    ,  -0.62            // 423
        ,  0.266    , -0.089            // 424
        ,  0.266    , -0.266            // 425
        ,  0.089    , -0.089            // 426
        ,  0.089    , -0.266            // 427
        ,  0.266    , -0.443            // 428
        ,  0.266    ,  -0.62            // 429
        ,  0.089    , -0.443            // 430
        ,  0.089    ,  -0.62            // 431
        ,   0.62    , -0.797            // 432
        ,   0.62    , -0.975            // 433
        ,  0.443    , -0.797            // 434
        ,  0.443    , -0.975            // 435
        ,   0.62    , -1.152            // 436
        ,   0.62    , -1.329            // 437
        ,  0.443    , -1.152            // 438
        ,  0.443    , -1.329            // 439
        ,  0.266    , -0.797            // 440
        ,  0.266    , -0.975            // 441
        ,  0.089    , -0.797            // 442
        ,  0.089    , -0.975            // 443
        ,  0.266    , -1.152            // 444
        ,  0.266    , -1.329            // 445
        ,  0.089    , -1.152            // 446
        ,  0.089    , -1.329            // 447
        ,  1.329    , -1.506            // 448
        ,  1.329    , -1.683            // 449
        ,  1.152    , -1.506            // 450
        ,  1.152    , -1.683            // 451
        ,  1.329    , -1.861            // 452
        ,  1.329    , -2.038            // 453
        ,  1.152    , -1.861            // 454
        ,  1.152    , -2.038            // 455
        ,  0.975    , -1.506            // 456
        ,  0.975    , -1.683            // 457
        ,  0.797    , -1.506            // 458
        ,  0.797    , -1.683            // 459
        ,  0.975    , -1.861            // 460
        ,  0.975    , -2.038            // 461
        ,  0.797    , -1.861            // 462
        ,  0.797    , -2.038            // 463
        ,  1.329    , -2.215            // 464
        ,  1.329    , -2.392            // 465
        ,  1.152    , -2.215            // 466
        ,  1.152    , -2.392            // 467
        ,  1.329    , -2.569            // 468
        ,  1.329    , -2.747            // 469
        ,  1.152    , -2.569            // 470
        ,  1.152    , -2.747            // 471
        ,  0.975    , -2.215            // 472
        ,  0.975    , -2.392            // 473
        ,  0.797    , -2.215            // 474
        ,  0.797    , -2.392            // 475
        ,  0.975    , -2.569            // 476
        ,  0.975    , -2.747            // 477
        ,  0.797    , -2.569            // 478
        ,  0.797    , -2.747            // 479
        ,   0.62    , -1.506            // 480
        ,   0.62    , -1.683            // 481
        ,  0.443    , -1.506            // 482
        ,  0.443    , -1.683            // 483
        ,   0.62    , -1.861            // 484
        ,   0.62    , -2.038            // 485
        ,  0.443    , -1.861            // 486
        ,  0.443    , -2.038            // 487
        ,  0.266    , -1.506            // 488
        ,  0.266    , -1.683            // 489
        ,  0.089    , -1.506            // 490
        ,  0.089    , -1.683            // 491
        ,  0.266    , -1.861            // 492
        ,  0.266    , -2.038            // 493
        ,  0.089    , -1.861            // 494
        ,  0.089    , -2.038            // 495
        ,   0.62    , -2.215            // 496
        ,   0.62    , -2.392            // 497
        ,  0.443    , -2.215            // 498
        ,  0.443    , -2.392            // 499
        ,   0.62    , -2.569            // 500
        ,   0.62    , -2.747            // 501
        ,  0.443    , -2.569            // 502
        ,  0.443    , -2.747            // 503
        ,  0.266    , -2.215            // 504
        ,  0.266    , -2.392            // 505
        ,  0.089    , -2.215            // 506
        ,  0.089    , -2.392            // 507
        ,  0.266    , -2.569            // 508
        ,  0.266    , -2.747            // 509
        ,  0.089    , -2.569            // 510
        ,  0.089    , -2.747            // 511
        , -0.089    ,  2.747            // 512
        , -0.089    ,  2.569            // 513
        , -0.266    ,  2.747            // 514
        , -0.266    ,  2.569            // 515
        , -0.089    ,  2.392            // 516
        , -0.089    ,  2.215            // 517
        , -0.266    ,  2.392            // 518
        , -0.266    ,  2.215            // 519
        , -0.443    ,  2.747            // 520
        , -0.443    ,  2.569            // 521
        ,  -0.62    ,  2.747            // 522
        ,  -0.62    ,  2.569            // 523
        , -0.443    ,  2.392            // 524
        , -0.443    ,  2.215            // 525
        ,  -0.62    ,  2.392            // 526
        ,  -0.62    ,  2.215            // 527
        , -0.089    ,  2.038            // 528
        , -0.089    ,  1.861            // 529
        , -0.266    ,  2.038            // 530
        , -0.266    ,  1.861            // 531
        , -0.089    ,  1.683            // 532
        , -0.089    ,  1.506            // 533
        , -0.266    ,  1.683            // 534
        , -0.266    ,  1.506            // 535
        , -0.443    ,  2.038            // 536
        , -0.443    ,  1.861            // 537
        ,  -0.62    ,  2.038            // 538
        ,  -0.62    ,  1.861            // 539
        , -0.443    ,  1.683            // 540
        , -0.443    ,  1.506            // 541
        ,  -0.62    ,  1.683            // 542
        ,  -0.62    ,  1.506            // 543
        , -0.797    ,  2.747            // 544
        , -0.797    ,  2.569            // 545
        , -0.975    ,  2.747            // 546
        , -0.975    ,  2.569            // 547
        , -0.797    ,  2.392            // 548
        , -0.797    ,  2.215            // 549
        , -0.975    ,  2.392            // 550
        , -0.975    ,  2.215            // 551
        , -1.152    ,  2.747            // 552
        , -1.152    ,  2.569            // 553
        , -1.329    ,  2.747            // 554
        , -1.329    ,  2.569            // 555
        , -1.152    ,  2.392            // 556
        , -1.152    ,  2.215            // 557
        , -1.329    ,  2.392            // 558
        , -1.329    ,  2.215            // 559
        , -0.797    ,  2.038            // 560
        , -0.797    ,  1.861            // 561
        , -0.975    ,  2.038            // 562
        , -0.975    ,  1.861            // 563
        , -0.797    ,  1.683            // 564
        , -0.797    ,  1.506            // 565
        , -0.975    ,  1.683            // 566
        , -0.975    ,  1.506            // 567
        , -1.152    ,  2.038            // 568
        , -1.152    ,  1.861            // 569
        , -1.329    ,  2.038            // 570
        , -1.329    ,  1.861            // 571
        , -1.152    ,  1.683            // 572
        , -1.152    ,  1.506            // 573
        , -1.329    ,  1.683            // 574
        , -1.329    ,  1.506            // 575
        , -0.089    ,  1.329            // 576
        , -0.089    ,  1.152            // 577
        , -0.266    ,  1.329            // 578
        , -0.266    ,  1.152            // 579
        , -0.089    ,  0.975            // 580
        , -0.089    ,  0.797            // 581
        , -0.266    ,  0.975            // 582
        , -0.266    ,  0.797            // 583
        , -0.443    ,  1.329            // 584
        , -0.443    ,  1.152            // 585
        ,  -0.62    ,  1.329            // 586
        ,  -0.62    ,  1.152            // 587
        , -0.443    ,  0.975            // 588
        , -0.443    ,  0.797            // 589
        ,  -0.62    ,  0.975            // 590
        ,  -0.62    ,  0.797            // 591
        , -0.089    ,   0.62            // 592
        , -0.089    ,  0.443            // 593
        , -0.266    ,   0.62            // 594
        , -0.266    ,  0.443            // 595
        , -0.089    ,  0.266            // 596
        , -0.089    ,  0.089            // 597
        , -0.266    ,  0.266            // 598
        , -0.266    ,  0.089            // 599
        , -0.443    ,   0.62            // 600
        , -0.443    ,  0.443            // 601
        ,  -0.62    ,   0.62            // 602
        ,  -0.62    ,  0.443            // 603
        , -0.443    ,  0.266            // 604
        , -0.443    ,  0.089            // 605
        ,  -0.62    ,  0.266            // 606
        ,  -0.62    ,  0.089            // 607
        , -0.797    ,  1.329            // 608
        , -0.797    ,  1.152            // 609
        , -0.975    ,  1.329            // 610
        , -0.975    ,  1.152            // 611
        , -0.797    ,  0.975            // 612
        , -0.797    ,  0.797            // 613
        , -0.975    ,  0.975            // 614
        , -0.975    ,  0.797            // 615
        , -1.152    ,  1.329            // 616
        , -1.152    ,  1.152            // 617
        , -1.329    ,  1.329            // 618
        , -1.329    ,  1.152            // 619
        , -1.152    ,  0.975            // 620
        , -1.152    ,  0.797            // 621
        , -1.329    ,  0.975            // 622
        , -1.329    ,  0.797            // 623
        , -0.797    ,   0.62            // 624
        , -0.797    ,  0.443            // 625
        , -0.975    ,   0.62            // 626
        , -0.975    ,  0.443            // 627
        , -0.797    ,  0.266            // 628
        , -0.797    ,  0.089            // 629
        , -0.975    ,  0.266            // 630
        , -0.975    ,  0.089            // 631
        , -1.152    ,   0.62            // 632
        , -1.152    ,  0.443            // 633
        , -1.329    ,   0.62            // 634
        , -1.329    ,  0.443            // 635
        , -1.152    ,  0.266            // 636
        , -1.152    ,  0.089            // 637
        , -1.329    ,  0.266            // 638
        , -1.329    ,  0.089            // 639
        , -1.506    ,  2.747            // 640
        , -1.506    ,  2.569            // 641
        , -1.683    ,  2.747            // 642
        , -1.683    ,  2.569            // 643
        , -1.506    ,  2.392            // 644
        , -1.506    ,  2.215            // 645
        , -1.683    ,  2.392            // 646
        , -1.683    ,  2.215            // 647
        , -1.861    ,  2.747            // 648
        , -1.861    ,  2.569            // 649
        , -2.038    ,  2.747            // 650
        , -2.038    ,  2.569            // 651
        , -1.861    ,  2.392            // 652
        , -1.861    ,  2.215            // 653
        , -2.038    ,  2.392            // 654
        , -2.038    ,  2.215            // 655
        , -1.506    ,  2.038            // 656
        , -1.506    ,  1.861            // 657
        , -1.683    ,  2.038            // 658
        , -1.683    ,  1.861            // 659
        , -1.506    ,  1.683            // 660
        , -1.506    ,  1.506            // 661
        , -1.683    ,  1.683            // 662
        , -1.683    ,  1.506            // 663
        , -1.861    ,  2.038            // 664
        , -1.861    ,  1.861            // 665
        , -2.038    ,  2.038            // 666
        , -2.038    ,  1.861            // 667
        , -1.861    ,  1.683            // 668
        , -1.861    ,  1.506            // 669
        , -2.038    ,  1.683            // 670
        , -2.038    ,  1.506            // 671
        , -2.215    ,  2.747            // 672
        , -2.215    ,  2.569            // 673
        , -2.392    ,  2.747            // 674
        , -2.392    ,  2.569            // 675
        , -2.215    ,  2.392            // 676
        , -2.215    ,  2.215            // 677
        , -2.392    ,  2.392            // 678
        , -2.392    ,  2.215            // 679
        , -2.569    ,  2.747            // 680
        , -2.569    ,  2.569            // 681
        , -2.747    ,  2.747            // 682
        , -2.747    ,  2.569            // 683
        , -2.569    ,  2.392            // 684
        , -2.569    ,  2.215            // 685
        , -2.747    ,  2.392            // 686
        , -2.747    ,  2.215            // 687
        , -2.215    ,  2.038            // 688
        , -2.215    ,  1.861            // 689
        , -2.392    ,  2.038            // 690
        , -2.392    ,  1.861            // 691
        , -2.215    ,  1.683            // 692
        , -2.215    ,  1.506            // 693
        , -2.392    ,  1.683            // 694
        , -2.392    ,  1.506            // 695
        , -2.569    ,  2.038            // 696
        , -2.569    ,  1.861            // 697
        , -2.747    ,  2.038            // 698
        , -2.747    ,  1.861            // 699
        , -2.569    ,  1.683            // 700
        , -2.569    ,  1.506            // 701
        , -2.747    ,  1.683            // 702
        , -2.747    ,  1.506            // 703
        , -1.506    ,  1.329            // 704
        , -1.506    ,  1.152            // 705
        , -1.683    ,  1.329            // 706
        , -1.683    ,  1.152            // 707
        , -1.506    ,  0.975            // 708
        , -1.506    ,  0.797            // 709
        , -1.683    ,  0.975            // 710
        , -1.683    ,  0.797            // 711
        , -1.861    ,  1.329            // 712
        , -1.861    ,  1.152            // 713
        , -2.038    ,  1.329            // 714
        , -2.038    ,  1.152            // 715
        , -1.861    ,  0.975            // 716
        , -1.861    ,  0.797            // 717
        , -2.038    ,  0.975            // 718
        , -2.038    ,  0.797            // 719
        , -1.506    ,   0.62            // 720
        , -1.506    ,  0.443            // 721
        , -1.683    ,   0.62            // 722
        , -1.683    ,  0.443            // 723
        , -1.506    ,  0.266            // 724
        , -1.506    ,  0.089            // 725
        , -1.683    ,  0.266            // 726
        , -1.683    ,  0.089            // 727
        , -1.861    ,   0.62            // 728
        , -1.861    ,  0.443            // 729
        , -2.038    ,   0.62            // 730
        , -2.038    ,  0.443            // 731
        , -1.861    ,  0.266            // 732
        , -1.861    ,  0.089            // 733
        , -2.038    ,  0.266            // 734
        , -2.038    ,  0.089            // 735
        , -2.215    ,  1.329            // 736
        , -2.215    ,  1.152            // 737
        , -2.392    ,  1.329            // 738
        , -2.392    ,  1.152            // 739
        , -2.215    ,  0.975            // 740
        , -2.215    ,  0.797            // 741
        , -2.392    ,  0.975            // 742
        , -2.392    ,  0.797            // 743
        , -2.569    ,  1.329            // 744
        , -2.569    ,  1.152            // 745
        , -2.747    ,  1.329            // 746
        , -2.747    ,  1.152            // 747
        , -2.569    ,  0.975            // 748
        , -2.569    ,  0.797            // 749
        , -2.747    ,  0.975            // 750
        , -2.747    ,  0.797            // 751
        , -2.215    ,   0.62            // 752
        , -2.215    ,  0.443            // 753
        , -2.392    ,   0.62            // 754
        , -2.392    ,  0.443            // 755
        , -2.215    ,  0.266            // 756
        , -2.215    ,  0.089            // 757
        , -2.392    ,  0.266            // 758
        , -2.392    ,  0.089            // 759
        , -2.569    ,   0.62            // 760
        , -2.569    ,  0.443            // 761
        , -2.747    ,   0.62            // 762
        , -2.747    ,  0.443            // 763
        , -2.569    ,  0.266            // 764
        , -2.569    ,  0.089            // 765
        , -2.747    ,  0.266            // 766
        , -2.747    ,  0.089            // 767
        , -0.089    , -0.089            // 768
        , -0.089    , -0.266            // 769
        , -0.266    , -0.089            // 770
        , -0.266    , -0.266            // 771
        , -0.089    , -0.443            // 772
        , -0.089    ,  -0.62            // 773
        , -0.266    , -0.443            // 774
        , -0.266    ,  -0.62            // 775
        , -0.443    , -0.089            // 776
        , -0.443    , -0.266            // 777
        ,  -0.62    , -0.089            // 778
        ,  -0.62    , -0.266            // 779
        , -0.443    , -0.443            // 780
        , -0.443    ,  -0.62            // 781
        ,  -0.62    , -0.443            // 782
        ,  -0.62    ,  -0.62            // 783
        , -0.089    , -0.797            // 784
        , -0.089    , -0.975            // 785
        , -0.266    , -0.797            // 786
        , -0.266    , -0.975            // 787
        , -0.089    , -1.152            // 788
        , -0.089    , -1.329            // 789
        , -0.266    , -1.152            // 790
        , -0.266    , -1.329            // 791
        , -0.443    , -0.797            // 792
        , -0.443    , -0.975            // 793
        ,  -0.62    , -0.797            // 794
        ,  -0.62    , -0.975            // 795
        , -0.443    , -1.152            // 796
        , -0.443    , -1.329            // 797
        ,  -0.62    , -1.152            // 798
        ,  -0.62    , -1.329            // 799
        , -0.797    , -0.089            // 800
        , -0.797    , -0.266            // 801
        , -0.975    , -0.089            // 802
        , -0.975    , -0.266            // 803
        , -0.797    , -0.443            // 804
        , -0.797    ,  -0.62            // 805
        , -0.975    , -0.443            // 806
        , -0.975    ,  -0.62            // 807
        , -1.152    , -0.089            // 808
        , -1.152    , -0.266            // 809
        , -1.329    , -0.089            // 810
        , -1.329    , -0.266            // 811
        , -1.152    , -0.443            // 812
        , -1.152    ,  -0.62            // 813
        , -1.329    , -0.443            // 814
        , -1.329    ,  -0.62            // 815
        , -0.797    , -0.797            // 816
        , -0.797    , -0.975            // 817
        , -0.975    , -0.797            // 818
        , -0.975    , -0.975            // 819
        , -0.797    , -1.152            // 820
        , -0.797    , -1.329            // 821
        , -0.975    , -1.152            // 822
        , -0.975    , -1.329            // 823
        , -1.152    , -0.797            // 824
        , -1.152    , -0.975            // 825
        , -1.329    , -0.797            // 826
        , -1.329    , -0.975            // 827
        , -1.152    , -1.152            // 828
        , -1.152    , -1.329            // 829
        , -1.329    , -1.152            // 830
        , -1.329    , -1.329            // 831
        , -0.089    , -1.506            // 832
        , -0.089    , -1.683            // 833
        , -0.266    , -1.506            // 834
        , -0.266    , -1.683            // 835
        , -0.089    , -1.861            // 836
        , -0.089    , -2.038            // 837
        , -0.266    , -1.861            // 838
        , -0.266    , -2.038            // 839
        , -0.443    , -1.506            // 840
        , -0.443    , -1.683            // 841
        ,  -0.62    , -1.506            // 842
        ,  -0.62    , -1.683            // 843
        , -0.443    , -1.861            // 844
        , -0.443    , -2.038            // 845
        ,  -0.62    , -1.861            // 846
        ,  -0.62    , -2.038            // 847
        , -0.089    , -2.215            // 848
        , -0.089    , -2.392            // 849
        , -0.266    , -2.215            // 850
        , -0.266    , -2.392            // 851
        , -0.089    , -2.569            // 852
        , -0.089    , -2.747            // 853
        , -0.266    , -2.569            // 854
        , -0.266    , -2.747            // 855
        , -0.443    , -2.215            // 856
        , -0.443    , -2.392            // 857
        ,  -0.62    , -2.215            // 858
        ,  -0.62    , -2.392            // 859
        , -0.443    , -2.569            // 860
        , -0.443    , -2.747            // 861
        ,  -0.62    , -2.569            // 862
        ,  -0.62    , -2.747            // 863
        , -0.797    , -1.506            // 864
        , -0.797    , -1.683            // 865
        , -0.975    , -1.506            // 866
        , -0.975    , -1.683            // 867
        , -0.797    , -1.861            // 868
        , -0.797    , -2.038            // 869
        , -0.975    , -1.861            // 870
        , -0.975    , -2.038            // 871
        , -1.152    , -1.506            // 872
        , -1.152    , -1.683            // 873
        , -1.329    , -1.506            // 874
        , -1.329    , -1.683            // 875
        , -1.152    , -1.861            // 876
        , -1.152    , -2.038            // 877
        , -1.329    , -1.861            // 878
        , -1.329    , -2.038            // 879
        , -0.797    , -2.215            // 880
        , -0.797    , -2.392            // 881
        , -0.975    , -2.215            // 882
        , -0.975    , -2.392            // 883
        , -0.797    , -2.569            // 884
        , -0.797    , -2.747            // 885
        , -0.975    , -2.569            // 886
        , -0.975    , -2.747            // 887
        , -1.152    , -2.215            // 888
        , -1.152    , -2.392            // 889
        , -1.329    , -2.215            // 890
        , -1.329    , -2.392            // 891
        , -1.152    , -2.569            // 892
        , -1.152    , -2.747            // 893
        , -1.329    , -2.569            // 894
        , -1.329    , -2.747            // 895
        , -1.506    , -0.089            // 896
        , -1.506    , -0.266            // 897
        , -1.683    , -0.089            // 898
        , -1.683    , -0.266            // 899
        , -1.506    , -0.443            // 900
        , -1.506    ,  -0.62            // 901
        , -1.683    , -0.443            // 902
        , -1.683    ,  -0.62            // 903
        , -1.861    , -0.089            // 904
        , -1.861    , -0.266            // 905
        , -2.038    , -0.089            // 906
        , -2.038    , -0.266            // 907
        , -1.861    , -0.443            // 908
        , -1.861    ,  -0.62            // 909
        , -2.038    , -0.443            // 910
        , -2.038    ,  -0.62            // 911
        , -1.506    , -0.797            // 912
        , -1.506    , -0.975            // 913
        , -1.683    , -0.797            // 914
        , -1.683    , -0.975            // 915
        , -1.506    , -1.152            // 916
        , -1.506    , -1.329            // 917
        , -1.683    , -1.152            // 918
        , -1.683    , -1.329            // 919
        , -1.861    , -0.797            // 920
        , -1.861    , -0.975            // 921
        , -2.038    , -0.797            // 922
        , -2.038    , -0.975            // 923
        , -1.861    , -1.152            // 924
        , -1.861    , -1.329            // 925
        , -2.038    , -1.152            // 926
        , -2.038    , -1.329            // 927
        , -2.215    , -0.089            // 928
        , -2.215    , -0.266            // 929
        , -2.392    , -0.089            // 930
        , -2.392    , -0.266            // 931
        , -2.215    , -0.443            // 932
        , -2.215    ,  -0.62            // 933
        , -2.392    , -0.443            // 934
        , -2.392    ,  -0.62            // 935
        , -2.569    , -0.089            // 936
        , -2.569    , -0.266            // 937
        , -2.747    , -0.089            // 938
        , -2.747    , -0.266            // 939
        , -2.569    , -0.443            // 940
        , -2.569    ,  -0.62            // 941
        , -2.747    , -0.443            // 942
        , -2.747    ,  -0.62            // 943
        , -2.215    , -0.797            // 944
        , -2.215    , -0.975            // 945
        , -2.392    , -0.797            // 946
        , -2.392    , -0.975            // 947
        , -2.215    , -1.152            // 948
        , -2.215    , -1.329            // 949
        , -2.392    , -1.152            // 950
        , -2.392    , -1.329            // 951
        , -2.569    , -0.797            // 952
        , -2.569    , -0.975            // 953
        , -2.747    , -0.797            // 954
        , -2.747    , -0.975            // 955
        , -2.569    , -1.152            // 956
        , -2.569    , -1.329            // 957
        , -2.747    , -1.152            // 958
        , -2.747    , -1.329            // 959
        , -1.506    , -1.506            // 960
        , -1.506    , -1.683            // 961
        , -1.683    , -1.506            // 962
        , -1.683    , -1.683            // 963
        , -1.506    , -1.861            // 964
        , -1.506    , -2.038            // 965
        , -1.683    , -1.861            // 966
        , -1.683    , -2.038            // 967
        , -1.861    , -1.506            // 968
        , -1.861    , -1.683            // 969
        , -2.038    , -1.506            // 970
        , -2.038    , -1.683            // 971
        , -1.861    , -1.861            // 972
        , -1.861    , -2.038            // 973
        , -2.038    , -1.861            // 974
        , -2.038    , -2.038            // 975
        , -1.506    , -2.215            // 976
        , -1.506    , -2.392            // 977
        , -1.683    , -2.215            // 978
        , -1.683    , -2.392            // 979
        , -1.506    , -2.569            // 980
        , -1.506    , -2.747            // 981
        , -1.683    , -2.569            // 982
        , -1.683    , -2.747            // 983
        , -1.861    , -2.215            // 984
        , -1.861    , -2.392            // 985
        , -2.038    , -2.215            // 986
        , -2.038    , -2.392            // 987
        , -1.861    , -2.569            // 988
        , -1.861    , -2.747            // 989
        , -2.038    , -2.569            // 990
        , -2.038    , -2.747            // 991
        , -2.215    , -1.506            // 992
        , -2.215    , -1.683            // 993
        , -2.392    , -1.506            // 994
        , -2.392    , -1.683            // 995
        , -2.215    , -1.861            // 996
        , -2.215    , -2.038            // 997
        , -2.392    , -1.861            // 998
        , -2.392    , -2.038            // 999
        , -2.569    , -1.506            // 1000
        , -2.569    , -1.683            // 1001
        , -2.747    , -1.506            // 1002
        , -2.747    , -1.683            // 1003
        , -2.569    , -1.861            // 1004
        , -2.569    , -2.038            // 1005
        , -2.747    , -1.861            // 1006
        , -2.747    , -2.038            // 1007
        , -2.215    , -2.215            // 1008
        , -2.215    , -2.392            // 1009
        , -2.392    , -2.215            // 1010
        , -2.392    , -2.392            // 1011
        , -2.215    , -2.569            // 1012
        , -2.215    , -2.747            // 1013
        , -2.392    , -2.569            // 1014
        , -2.392    , -2.747            // 1015
        , -2.569    , -2.215            // 1016
        , -2.569    , -2.392            // 1017
        , -2.747    , -2.215            // 1018
        , -2.747    , -2.392            // 1019
        , -2.569    , -2.569            // 1020
        , -2.569    , -2.747            // 1021
        , -2.747    , -2.569            // 1022
        , -2.747    , -2.747            // 1023
    };