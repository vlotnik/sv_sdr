    DVBS2X_8_16_20_20APSK_5_6 : super.plane = {
           0.119    , -0.599            // 0
        ,  0.981    , -0.981            // 1
        ,  0.339    , -0.508            // 2
        ,  0.687    , -0.687            // 3
        ,  0.217    , -1.371            // 4
        ,   0.63    , -1.237            // 5
        ,  0.152    ,  -0.96            // 6
        ,  0.441    , -0.866            // 7
        , -0.119    , -0.599            // 8
        , -0.981    , -0.981            // 9
        , -0.339    , -0.508            // 10
        , -0.687    , -0.687            // 11
        , -0.217    , -1.371            // 12
        ,  -0.63    , -1.237            // 13
        , -0.152    ,  -0.96            // 14
        , -0.441    , -0.866            // 15
        ,  0.106    , -0.256            // 16
        ,  1.237    ,  -0.63            // 17
        ,  0.508    , -0.339            // 18
        ,  0.866    , -0.441            // 19
        ,  0.256    , -0.106            // 20
        ,  1.371    , -0.217            // 21
        ,  0.599    , -0.119            // 22
        ,   0.96    , -0.152            // 23
        , -0.106    , -0.256            // 24
        , -1.237    ,  -0.63            // 25
        , -0.508    , -0.339            // 26
        , -0.866    , -0.441            // 27
        , -0.256    , -0.106            // 28
        , -1.371    , -0.217            // 29
        , -0.599    , -0.119            // 30
        ,  -0.96    , -0.152            // 31
        ,  0.119    ,  0.599            // 32
        ,  0.981    ,  0.981            // 33
        ,  0.339    ,  0.508            // 34
        ,  0.687    ,  0.687            // 35
        ,  0.217    ,  1.371            // 36
        ,   0.63    ,  1.237            // 37
        ,  0.152    ,   0.96            // 38
        ,  0.441    ,  0.866            // 39
        , -0.119    ,  0.599            // 40
        , -0.981    ,  0.981            // 41
        , -0.339    ,  0.508            // 42
        , -0.687    ,  0.687            // 43
        , -0.217    ,  1.371            // 44
        ,  -0.63    ,  1.237            // 45
        , -0.152    ,   0.96            // 46
        , -0.441    ,  0.866            // 47
        ,  0.106    ,  0.256            // 48
        ,  1.237    ,   0.63            // 49
        ,  0.508    ,  0.339            // 50
        ,  0.866    ,  0.441            // 51
        ,  0.256    ,  0.106            // 52
        ,  1.371    ,  0.217            // 53
        ,  0.599    ,  0.119            // 54
        ,   0.96    ,  0.152            // 55
        , -0.106    ,  0.256            // 56
        , -1.237    ,   0.63            // 57
        , -0.508    ,  0.339            // 58
        , -0.866    ,  0.441            // 59
        , -0.256    ,  0.106            // 60
        , -1.371    ,  0.217            // 61
        , -0.599    ,  0.119            // 62
        ,  -0.96    ,  0.152            // 63
    };