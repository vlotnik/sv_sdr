    QAM256 : super.plane = {
           1.335    ,  1.335            // 0
        ,  1.335    ,  1.157            // 1
        ,  1.157    ,  1.335            // 2
        ,  1.157    ,  1.157            // 3
        ,  1.335    ,  0.979            // 4
        ,  1.335    ,  0.801            // 5
        ,  1.157    ,  0.979            // 6
        ,  1.157    ,  0.801            // 7
        ,  0.979    ,  1.335            // 8
        ,  0.979    ,  1.157            // 9
        ,  0.801    ,  1.335            // 10
        ,  0.801    ,  1.157            // 11
        ,  0.979    ,  0.979            // 12
        ,  0.979    ,  0.801            // 13
        ,  0.801    ,  0.979            // 14
        ,  0.801    ,  0.801            // 15
        ,  1.335    ,  0.623            // 16
        ,  1.335    ,  0.445            // 17
        ,  1.157    ,  0.623            // 18
        ,  1.157    ,  0.445            // 19
        ,  1.335    ,  0.267            // 20
        ,  1.335    ,  0.089            // 21
        ,  1.157    ,  0.267            // 22
        ,  1.157    ,  0.089            // 23
        ,  0.979    ,  0.623            // 24
        ,  0.979    ,  0.445            // 25
        ,  0.801    ,  0.623            // 26
        ,  0.801    ,  0.445            // 27
        ,  0.979    ,  0.267            // 28
        ,  0.979    ,  0.089            // 29
        ,  0.801    ,  0.267            // 30
        ,  0.801    ,  0.089            // 31
        ,  0.623    ,  1.335            // 32
        ,  0.623    ,  1.157            // 33
        ,  0.445    ,  1.335            // 34
        ,  0.445    ,  1.157            // 35
        ,  0.623    ,  0.979            // 36
        ,  0.623    ,  0.801            // 37
        ,  0.445    ,  0.979            // 38
        ,  0.445    ,  0.801            // 39
        ,  0.267    ,  1.335            // 40
        ,  0.267    ,  1.157            // 41
        ,  0.089    ,  1.335            // 42
        ,  0.089    ,  1.157            // 43
        ,  0.267    ,  0.979            // 44
        ,  0.267    ,  0.801            // 45
        ,  0.089    ,  0.979            // 46
        ,  0.089    ,  0.801            // 47
        ,  0.623    ,  0.623            // 48
        ,  0.623    ,  0.445            // 49
        ,  0.445    ,  0.623            // 50
        ,  0.445    ,  0.445            // 51
        ,  0.623    ,  0.267            // 52
        ,  0.623    ,  0.089            // 53
        ,  0.445    ,  0.267            // 54
        ,  0.445    ,  0.089            // 55
        ,  0.267    ,  0.623            // 56
        ,  0.267    ,  0.445            // 57
        ,  0.089    ,  0.623            // 58
        ,  0.089    ,  0.445            // 59
        ,  0.267    ,  0.267            // 60
        ,  0.267    ,  0.089            // 61
        ,  0.089    ,  0.267            // 62
        ,  0.089    ,  0.089            // 63
        ,  1.335    , -0.089            // 64
        ,  1.335    , -0.267            // 65
        ,  1.157    , -0.089            // 66
        ,  1.157    , -0.267            // 67
        ,  1.335    , -0.445            // 68
        ,  1.335    , -0.623            // 69
        ,  1.157    , -0.445            // 70
        ,  1.157    , -0.623            // 71
        ,  0.979    , -0.089            // 72
        ,  0.979    , -0.267            // 73
        ,  0.801    , -0.089            // 74
        ,  0.801    , -0.267            // 75
        ,  0.979    , -0.445            // 76
        ,  0.979    , -0.623            // 77
        ,  0.801    , -0.445            // 78
        ,  0.801    , -0.623            // 79
        ,  1.335    , -0.801            // 80
        ,  1.335    , -0.979            // 81
        ,  1.157    , -0.801            // 82
        ,  1.157    , -0.979            // 83
        ,  1.335    , -1.157            // 84
        ,  1.335    , -1.335            // 85
        ,  1.157    , -1.157            // 86
        ,  1.157    , -1.335            // 87
        ,  0.979    , -0.801            // 88
        ,  0.979    , -0.979            // 89
        ,  0.801    , -0.801            // 90
        ,  0.801    , -0.979            // 91
        ,  0.979    , -1.157            // 92
        ,  0.979    , -1.335            // 93
        ,  0.801    , -1.157            // 94
        ,  0.801    , -1.335            // 95
        ,  0.623    , -0.089            // 96
        ,  0.623    , -0.267            // 97
        ,  0.445    , -0.089            // 98
        ,  0.445    , -0.267            // 99
        ,  0.623    , -0.445            // 100
        ,  0.623    , -0.623            // 101
        ,  0.445    , -0.445            // 102
        ,  0.445    , -0.623            // 103
        ,  0.267    , -0.089            // 104
        ,  0.267    , -0.267            // 105
        ,  0.089    , -0.089            // 106
        ,  0.089    , -0.267            // 107
        ,  0.267    , -0.445            // 108
        ,  0.267    , -0.623            // 109
        ,  0.089    , -0.445            // 110
        ,  0.089    , -0.623            // 111
        ,  0.623    , -0.801            // 112
        ,  0.623    , -0.979            // 113
        ,  0.445    , -0.801            // 114
        ,  0.445    , -0.979            // 115
        ,  0.623    , -1.157            // 116
        ,  0.623    , -1.335            // 117
        ,  0.445    , -1.157            // 118
        ,  0.445    , -1.335            // 119
        ,  0.267    , -0.801            // 120
        ,  0.267    , -0.979            // 121
        ,  0.089    , -0.801            // 122
        ,  0.089    , -0.979            // 123
        ,  0.267    , -1.157            // 124
        ,  0.267    , -1.335            // 125
        ,  0.089    , -1.157            // 126
        ,  0.089    , -1.335            // 127
        , -0.089    ,  1.335            // 128
        , -0.089    ,  1.157            // 129
        , -0.267    ,  1.335            // 130
        , -0.267    ,  1.157            // 131
        , -0.089    ,  0.979            // 132
        , -0.089    ,  0.801            // 133
        , -0.267    ,  0.979            // 134
        , -0.267    ,  0.801            // 135
        , -0.445    ,  1.335            // 136
        , -0.445    ,  1.157            // 137
        , -0.623    ,  1.335            // 138
        , -0.623    ,  1.157            // 139
        , -0.445    ,  0.979            // 140
        , -0.445    ,  0.801            // 141
        , -0.623    ,  0.979            // 142
        , -0.623    ,  0.801            // 143
        , -0.089    ,  0.623            // 144
        , -0.089    ,  0.445            // 145
        , -0.267    ,  0.623            // 146
        , -0.267    ,  0.445            // 147
        , -0.089    ,  0.267            // 148
        , -0.089    ,  0.089            // 149
        , -0.267    ,  0.267            // 150
        , -0.267    ,  0.089            // 151
        , -0.445    ,  0.623            // 152
        , -0.445    ,  0.445            // 153
        , -0.623    ,  0.623            // 154
        , -0.623    ,  0.445            // 155
        , -0.445    ,  0.267            // 156
        , -0.445    ,  0.089            // 157
        , -0.623    ,  0.267            // 158
        , -0.623    ,  0.089            // 159
        , -0.801    ,  1.335            // 160
        , -0.801    ,  1.157            // 161
        , -0.979    ,  1.335            // 162
        , -0.979    ,  1.157            // 163
        , -0.801    ,  0.979            // 164
        , -0.801    ,  0.801            // 165
        , -0.979    ,  0.979            // 166
        , -0.979    ,  0.801            // 167
        , -1.157    ,  1.335            // 168
        , -1.157    ,  1.157            // 169
        , -1.335    ,  1.335            // 170
        , -1.335    ,  1.157            // 171
        , -1.157    ,  0.979            // 172
        , -1.157    ,  0.801            // 173
        , -1.335    ,  0.979            // 174
        , -1.335    ,  0.801            // 175
        , -0.801    ,  0.623            // 176
        , -0.801    ,  0.445            // 177
        , -0.979    ,  0.623            // 178
        , -0.979    ,  0.445            // 179
        , -0.801    ,  0.267            // 180
        , -0.801    ,  0.089            // 181
        , -0.979    ,  0.267            // 182
        , -0.979    ,  0.089            // 183
        , -1.157    ,  0.623            // 184
        , -1.157    ,  0.445            // 185
        , -1.335    ,  0.623            // 186
        , -1.335    ,  0.445            // 187
        , -1.157    ,  0.267            // 188
        , -1.157    ,  0.089            // 189
        , -1.335    ,  0.267            // 190
        , -1.335    ,  0.089            // 191
        , -0.089    , -0.089            // 192
        , -0.089    , -0.267            // 193
        , -0.267    , -0.089            // 194
        , -0.267    , -0.267            // 195
        , -0.089    , -0.445            // 196
        , -0.089    , -0.623            // 197
        , -0.267    , -0.445            // 198
        , -0.267    , -0.623            // 199
        , -0.445    , -0.089            // 200
        , -0.445    , -0.267            // 201
        , -0.623    , -0.089            // 202
        , -0.623    , -0.267            // 203
        , -0.445    , -0.445            // 204
        , -0.445    , -0.623            // 205
        , -0.623    , -0.445            // 206
        , -0.623    , -0.623            // 207
        , -0.089    , -0.801            // 208
        , -0.089    , -0.979            // 209
        , -0.267    , -0.801            // 210
        , -0.267    , -0.979            // 211
        , -0.089    , -1.157            // 212
        , -0.089    , -1.335            // 213
        , -0.267    , -1.157            // 214
        , -0.267    , -1.335            // 215
        , -0.445    , -0.801            // 216
        , -0.445    , -0.979            // 217
        , -0.623    , -0.801            // 218
        , -0.623    , -0.979            // 219
        , -0.445    , -1.157            // 220
        , -0.445    , -1.335            // 221
        , -0.623    , -1.157            // 222
        , -0.623    , -1.335            // 223
        , -0.801    , -0.089            // 224
        , -0.801    , -0.267            // 225
        , -0.979    , -0.089            // 226
        , -0.979    , -0.267            // 227
        , -0.801    , -0.445            // 228
        , -0.801    , -0.623            // 229
        , -0.979    , -0.445            // 230
        , -0.979    , -0.623            // 231
        , -1.157    , -0.089            // 232
        , -1.157    , -0.267            // 233
        , -1.335    , -0.089            // 234
        , -1.335    , -0.267            // 235
        , -1.157    , -0.445            // 236
        , -1.157    , -0.623            // 237
        , -1.335    , -0.445            // 238
        , -1.335    , -0.623            // 239
        , -0.801    , -0.801            // 240
        , -0.801    , -0.979            // 241
        , -0.979    , -0.801            // 242
        , -0.979    , -0.979            // 243
        , -0.801    , -1.157            // 244
        , -0.801    , -1.335            // 245
        , -0.979    , -1.157            // 246
        , -0.979    , -1.335            // 247
        , -1.157    , -0.801            // 248
        , -1.157    , -0.979            // 249
        , -1.335    , -0.801            // 250
        , -1.335    , -0.979            // 251
        , -1.157    , -1.157            // 252
        , -1.157    , -1.335            // 253
        , -1.335    , -1.157            // 254
        , -1.335    , -1.335            // 255
    };