    DVBS2X_4_8_4_16APSK_140_180 : super.plane = {
           0.162    ,  0.162            // 0
        ,  0.251    ,  1.262            // 1
        ,  0.162    , -0.162            // 2
        ,  0.251    , -1.262            // 3
        , -0.162    ,  0.162            // 4
        , -0.251    ,  1.262            // 5
        , -0.162    , -0.162            // 6
        , -0.251    , -1.262            // 7
        ,  0.621    ,  0.166            // 8
        ,  1.262    ,  0.251            // 9
        ,  0.621    , -0.166            // 10
        ,  1.262    , -0.251            // 11
        , -0.621    ,  0.166            // 12
        , -1.262    ,  0.251            // 13
        , -0.621    , -0.166            // 14
        , -1.262    , -0.251            // 15
        ,  0.166    ,  0.621            // 16
        ,  0.715    ,   1.07            // 17
        ,  0.166    , -0.621            // 18
        ,  0.715    ,  -1.07            // 19
        , -0.166    ,  0.621            // 20
        , -0.715    ,   1.07            // 21
        , -0.166    , -0.621            // 22
        , -0.715    ,  -1.07            // 23
        ,    0.5    ,    0.5            // 24
        ,   1.07    ,  0.715            // 25
        ,    0.5    ,   -0.5            // 26
        ,   1.07    , -0.715            // 27
        ,   -0.5    ,    0.5            // 28
        ,  -1.07    ,  0.715            // 29
        ,   -0.5    ,   -0.5            // 30
        ,  -1.07    , -0.715            // 31
    };