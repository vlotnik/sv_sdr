    DVBS2_APSK32_5_6 : super.plane = {
           0.508    ,  0.508            // 0
        ,  0.186    ,  0.694            // 1
        ,  0.508    , -0.508            // 2
        ,  0.186    , -0.694            // 3
        , -0.508    ,  0.508            // 4
        , -0.186    ,  0.694            // 5
        , -0.508    , -0.508            // 6
        , -0.186    , -0.694            // 7
        ,  1.167    ,  0.483            // 8
        ,  0.483    ,  1.167            // 9
        ,  0.893    , -0.893            // 10
        ,      0    , -1.263            // 11
        , -0.893    ,  0.893            // 12
        ,      0    ,  1.263            // 13
        , -1.167    , -0.483            // 14
        , -0.483    , -1.167            // 15
        ,  0.694    ,  0.186            // 16
        ,  0.192    ,  0.192            // 17
        ,  0.694    , -0.186            // 18
        ,  0.192    , -0.192            // 19
        , -0.694    ,  0.186            // 20
        , -0.192    ,  0.192            // 21
        , -0.694    , -0.186            // 22
        , -0.192    , -0.192            // 23
        ,  1.263    ,      0            // 24
        ,  0.893    ,  0.893            // 25
        ,  1.167    , -0.483            // 26
        ,  0.483    , -1.167            // 27
        , -1.167    ,  0.483            // 28
        , -0.483    ,  1.167            // 29
        , -1.263    ,      0            // 30
        , -0.893    , -0.893            // 31
    };