    QAM512 : super.plane = {
           2.024    ,   1.32            // 0
        ,  2.024    ,  1.144            // 1
        ,  1.848    ,   1.32            // 2
        ,  1.848    ,  1.144            // 3
        ,  2.024    ,  0.968            // 4
        ,  2.024    ,  0.792            // 5
        ,  1.848    ,  0.968            // 6
        ,  1.848    ,  0.792            // 7
        ,  1.672    ,   1.32            // 8
        ,  1.672    ,  1.144            // 9
        ,  1.496    ,   1.32            // 10
        ,  1.496    ,  1.144            // 11
        ,  1.672    ,  0.968            // 12
        ,  1.672    ,  0.792            // 13
        ,  1.496    ,  0.968            // 14
        ,  1.496    ,  0.792            // 15
        ,  2.024    ,  0.616            // 16
        ,  2.024    ,   0.44            // 17
        ,  1.848    ,  0.616            // 18
        ,  1.848    ,   0.44            // 19
        ,  2.024    ,  0.264            // 20
        ,  2.024    ,  0.088            // 21
        ,  1.848    ,  0.264            // 22
        ,  1.848    ,  0.088            // 23
        ,  1.672    ,  0.616            // 24
        ,  1.672    ,   0.44            // 25
        ,  1.496    ,  0.616            // 26
        ,  1.496    ,   0.44            // 27
        ,  1.672    ,  0.264            // 28
        ,  1.672    ,  0.088            // 29
        ,  1.496    ,  0.264            // 30
        ,  1.496    ,  0.088            // 31
        ,   1.32    ,  2.024            // 32
        ,   1.32    ,  1.848            // 33
        ,  1.144    ,  2.024            // 34
        ,  1.144    ,  1.848            // 35
        ,   1.32    ,  1.672            // 36
        ,   1.32    ,  1.496            // 37
        ,  1.144    ,  1.672            // 38
        ,  1.144    ,  1.496            // 39
        ,  0.968    ,  2.024            // 40
        ,  0.968    ,  1.848            // 41
        ,  0.792    ,  2.024            // 42
        ,  0.792    ,  1.848            // 43
        ,  0.968    ,  1.672            // 44
        ,  0.968    ,  1.496            // 45
        ,  0.792    ,  1.672            // 46
        ,  0.792    ,  1.496            // 47
        ,  0.616    ,  2.024            // 48
        ,  0.616    ,  1.848            // 49
        ,   0.44    ,  2.024            // 50
        ,   0.44    ,  1.848            // 51
        ,  0.616    ,  1.672            // 52
        ,  0.616    ,  1.496            // 53
        ,   0.44    ,  1.672            // 54
        ,   0.44    ,  1.496            // 55
        ,  0.264    ,  2.024            // 56
        ,  0.264    ,  1.848            // 57
        ,  0.088    ,  2.024            // 58
        ,  0.088    ,  1.848            // 59
        ,  0.264    ,  1.672            // 60
        ,  0.264    ,  1.496            // 61
        ,  0.088    ,  1.672            // 62
        ,  0.088    ,  1.496            // 63
        ,   1.32    ,   1.32            // 64
        ,   1.32    ,  1.144            // 65
        ,  1.144    ,   1.32            // 66
        ,  1.144    ,  1.144            // 67
        ,   1.32    ,  0.968            // 68
        ,   1.32    ,  0.792            // 69
        ,  1.144    ,  0.968            // 70
        ,  1.144    ,  0.792            // 71
        ,  0.968    ,   1.32            // 72
        ,  0.968    ,  1.144            // 73
        ,  0.792    ,   1.32            // 74
        ,  0.792    ,  1.144            // 75
        ,  0.968    ,  0.968            // 76
        ,  0.968    ,  0.792            // 77
        ,  0.792    ,  0.968            // 78
        ,  0.792    ,  0.792            // 79
        ,   1.32    ,  0.616            // 80
        ,   1.32    ,   0.44            // 81
        ,  1.144    ,  0.616            // 82
        ,  1.144    ,   0.44            // 83
        ,   1.32    ,  0.264            // 84
        ,   1.32    ,  0.088            // 85
        ,  1.144    ,  0.264            // 86
        ,  1.144    ,  0.088            // 87
        ,  0.968    ,  0.616            // 88
        ,  0.968    ,   0.44            // 89
        ,  0.792    ,  0.616            // 90
        ,  0.792    ,   0.44            // 91
        ,  0.968    ,  0.264            // 92
        ,  0.968    ,  0.088            // 93
        ,  0.792    ,  0.264            // 94
        ,  0.792    ,  0.088            // 95
        ,  0.616    ,   1.32            // 96
        ,  0.616    ,  1.144            // 97
        ,   0.44    ,   1.32            // 98
        ,   0.44    ,  1.144            // 99
        ,  0.616    ,  0.968            // 100
        ,  0.616    ,  0.792            // 101
        ,   0.44    ,  0.968            // 102
        ,   0.44    ,  0.792            // 103
        ,  0.264    ,   1.32            // 104
        ,  0.264    ,  1.144            // 105
        ,  0.088    ,   1.32            // 106
        ,  0.088    ,  1.144            // 107
        ,  0.264    ,  0.968            // 108
        ,  0.264    ,  0.792            // 109
        ,  0.088    ,  0.968            // 110
        ,  0.088    ,  0.792            // 111
        ,  0.616    ,  0.616            // 112
        ,  0.616    ,   0.44            // 113
        ,   0.44    ,  0.616            // 114
        ,   0.44    ,   0.44            // 115
        ,  0.616    ,  0.264            // 116
        ,  0.616    ,  0.088            // 117
        ,   0.44    ,  0.264            // 118
        ,   0.44    ,  0.088            // 119
        ,  0.264    ,  0.616            // 120
        ,  0.264    ,   0.44            // 121
        ,  0.088    ,  0.616            // 122
        ,  0.088    ,   0.44            // 123
        ,  0.264    ,  0.264            // 124
        ,  0.264    ,  0.088            // 125
        ,  0.088    ,  0.264            // 126
        ,  0.088    ,  0.088            // 127
        ,  2.024    , -0.088            // 128
        ,  2.024    , -0.264            // 129
        ,  1.848    , -0.088            // 130
        ,  1.848    , -0.264            // 131
        ,  2.024    ,  -0.44            // 132
        ,  2.024    , -0.616            // 133
        ,  1.848    ,  -0.44            // 134
        ,  1.848    , -0.616            // 135
        ,  1.672    , -0.088            // 136
        ,  1.672    , -0.264            // 137
        ,  1.496    , -0.088            // 138
        ,  1.496    , -0.264            // 139
        ,  1.672    ,  -0.44            // 140
        ,  1.672    , -0.616            // 141
        ,  1.496    ,  -0.44            // 142
        ,  1.496    , -0.616            // 143
        ,  2.024    , -0.792            // 144
        ,  2.024    , -0.968            // 145
        ,  1.848    , -0.792            // 146
        ,  1.848    , -0.968            // 147
        ,  2.024    , -1.144            // 148
        ,  2.024    ,  -1.32            // 149
        ,  1.848    , -1.144            // 150
        ,  1.848    ,  -1.32            // 151
        ,  1.672    , -0.792            // 152
        ,  1.672    , -0.968            // 153
        ,  1.496    , -0.792            // 154
        ,  1.496    , -0.968            // 155
        ,  1.672    , -1.144            // 156
        ,  1.672    ,  -1.32            // 157
        ,  1.496    , -1.144            // 158
        ,  1.496    ,  -1.32            // 159
        ,   1.32    , -0.088            // 160
        ,   1.32    , -0.264            // 161
        ,  1.144    , -0.088            // 162
        ,  1.144    , -0.264            // 163
        ,   1.32    ,  -0.44            // 164
        ,   1.32    , -0.616            // 165
        ,  1.144    ,  -0.44            // 166
        ,  1.144    , -0.616            // 167
        ,  0.968    , -0.088            // 168
        ,  0.968    , -0.264            // 169
        ,  0.792    , -0.088            // 170
        ,  0.792    , -0.264            // 171
        ,  0.968    ,  -0.44            // 172
        ,  0.968    , -0.616            // 173
        ,  0.792    ,  -0.44            // 174
        ,  0.792    , -0.616            // 175
        ,   1.32    , -0.792            // 176
        ,   1.32    , -0.968            // 177
        ,  1.144    , -0.792            // 178
        ,  1.144    , -0.968            // 179
        ,   1.32    , -1.144            // 180
        ,   1.32    ,  -1.32            // 181
        ,  1.144    , -1.144            // 182
        ,  1.144    ,  -1.32            // 183
        ,  0.968    , -0.792            // 184
        ,  0.968    , -0.968            // 185
        ,  0.792    , -0.792            // 186
        ,  0.792    , -0.968            // 187
        ,  0.968    , -1.144            // 188
        ,  0.968    ,  -1.32            // 189
        ,  0.792    , -1.144            // 190
        ,  0.792    ,  -1.32            // 191
        ,  0.616    , -0.088            // 192
        ,  0.616    , -0.264            // 193
        ,   0.44    , -0.088            // 194
        ,   0.44    , -0.264            // 195
        ,  0.616    ,  -0.44            // 196
        ,  0.616    , -0.616            // 197
        ,   0.44    ,  -0.44            // 198
        ,   0.44    , -0.616            // 199
        ,  0.264    , -0.088            // 200
        ,  0.264    , -0.264            // 201
        ,  0.088    , -0.088            // 202
        ,  0.088    , -0.264            // 203
        ,  0.264    ,  -0.44            // 204
        ,  0.264    , -0.616            // 205
        ,  0.088    ,  -0.44            // 206
        ,  0.088    , -0.616            // 207
        ,  0.616    , -0.792            // 208
        ,  0.616    , -0.968            // 209
        ,   0.44    , -0.792            // 210
        ,   0.44    , -0.968            // 211
        ,  0.616    , -1.144            // 212
        ,  0.616    ,  -1.32            // 213
        ,   0.44    , -1.144            // 214
        ,   0.44    ,  -1.32            // 215
        ,  0.264    , -0.792            // 216
        ,  0.264    , -0.968            // 217
        ,  0.088    , -0.792            // 218
        ,  0.088    , -0.968            // 219
        ,  0.264    , -1.144            // 220
        ,  0.264    ,  -1.32            // 221
        ,  0.088    , -1.144            // 222
        ,  0.088    ,  -1.32            // 223
        ,   1.32    , -1.496            // 224
        ,   1.32    , -1.672            // 225
        ,  1.144    , -1.496            // 226
        ,  1.144    , -1.672            // 227
        ,   1.32    , -1.848            // 228
        ,   1.32    , -2.024            // 229
        ,  1.144    , -1.848            // 230
        ,  1.144    , -2.024            // 231
        ,  0.968    , -1.496            // 232
        ,  0.968    , -1.672            // 233
        ,  0.792    , -1.496            // 234
        ,  0.792    , -1.672            // 235
        ,  0.968    , -1.848            // 236
        ,  0.968    , -2.024            // 237
        ,  0.792    , -1.848            // 238
        ,  0.792    , -2.024            // 239
        ,  0.616    , -1.496            // 240
        ,  0.616    , -1.672            // 241
        ,   0.44    , -1.496            // 242
        ,   0.44    , -1.672            // 243
        ,  0.616    , -1.848            // 244
        ,  0.616    , -2.024            // 245
        ,   0.44    , -1.848            // 246
        ,   0.44    , -2.024            // 247
        ,  0.264    , -1.496            // 248
        ,  0.264    , -1.672            // 249
        ,  0.088    , -1.496            // 250
        ,  0.088    , -1.672            // 251
        ,  0.264    , -1.848            // 252
        ,  0.264    , -2.024            // 253
        ,  0.088    , -1.848            // 254
        ,  0.088    , -2.024            // 255
        , -0.088    ,  2.024            // 256
        , -0.088    ,  1.848            // 257
        , -0.264    ,  2.024            // 258
        , -0.264    ,  1.848            // 259
        , -0.088    ,  1.672            // 260
        , -0.088    ,  1.496            // 261
        , -0.264    ,  1.672            // 262
        , -0.264    ,  1.496            // 263
        ,  -0.44    ,  2.024            // 264
        ,  -0.44    ,  1.848            // 265
        , -0.616    ,  2.024            // 266
        , -0.616    ,  1.848            // 267
        ,  -0.44    ,  1.672            // 268
        ,  -0.44    ,  1.496            // 269
        , -0.616    ,  1.672            // 270
        , -0.616    ,  1.496            // 271
        , -0.792    ,  2.024            // 272
        , -0.792    ,  1.848            // 273
        , -0.968    ,  2.024            // 274
        , -0.968    ,  1.848            // 275
        , -0.792    ,  1.672            // 276
        , -0.792    ,  1.496            // 277
        , -0.968    ,  1.672            // 278
        , -0.968    ,  1.496            // 279
        , -1.144    ,  2.024            // 280
        , -1.144    ,  1.848            // 281
        ,  -1.32    ,  2.024            // 282
        ,  -1.32    ,  1.848            // 283
        , -1.144    ,  1.672            // 284
        , -1.144    ,  1.496            // 285
        ,  -1.32    ,  1.672            // 286
        ,  -1.32    ,  1.496            // 287
        , -0.088    ,   1.32            // 288
        , -0.088    ,  1.144            // 289
        , -0.264    ,   1.32            // 290
        , -0.264    ,  1.144            // 291
        , -0.088    ,  0.968            // 292
        , -0.088    ,  0.792            // 293
        , -0.264    ,  0.968            // 294
        , -0.264    ,  0.792            // 295
        ,  -0.44    ,   1.32            // 296
        ,  -0.44    ,  1.144            // 297
        , -0.616    ,   1.32            // 298
        , -0.616    ,  1.144            // 299
        ,  -0.44    ,  0.968            // 300
        ,  -0.44    ,  0.792            // 301
        , -0.616    ,  0.968            // 302
        , -0.616    ,  0.792            // 303
        , -0.088    ,  0.616            // 304
        , -0.088    ,   0.44            // 305
        , -0.264    ,  0.616            // 306
        , -0.264    ,   0.44            // 307
        , -0.088    ,  0.264            // 308
        , -0.088    ,  0.088            // 309
        , -0.264    ,  0.264            // 310
        , -0.264    ,  0.088            // 311
        ,  -0.44    ,  0.616            // 312
        ,  -0.44    ,   0.44            // 313
        , -0.616    ,  0.616            // 314
        , -0.616    ,   0.44            // 315
        ,  -0.44    ,  0.264            // 316
        ,  -0.44    ,  0.088            // 317
        , -0.616    ,  0.264            // 318
        , -0.616    ,  0.088            // 319
        , -0.792    ,   1.32            // 320
        , -0.792    ,  1.144            // 321
        , -0.968    ,   1.32            // 322
        , -0.968    ,  1.144            // 323
        , -0.792    ,  0.968            // 324
        , -0.792    ,  0.792            // 325
        , -0.968    ,  0.968            // 326
        , -0.968    ,  0.792            // 327
        , -1.144    ,   1.32            // 328
        , -1.144    ,  1.144            // 329
        ,  -1.32    ,   1.32            // 330
        ,  -1.32    ,  1.144            // 331
        , -1.144    ,  0.968            // 332
        , -1.144    ,  0.792            // 333
        ,  -1.32    ,  0.968            // 334
        ,  -1.32    ,  0.792            // 335
        , -0.792    ,  0.616            // 336
        , -0.792    ,   0.44            // 337
        , -0.968    ,  0.616            // 338
        , -0.968    ,   0.44            // 339
        , -0.792    ,  0.264            // 340
        , -0.792    ,  0.088            // 341
        , -0.968    ,  0.264            // 342
        , -0.968    ,  0.088            // 343
        , -1.144    ,  0.616            // 344
        , -1.144    ,   0.44            // 345
        ,  -1.32    ,  0.616            // 346
        ,  -1.32    ,   0.44            // 347
        , -1.144    ,  0.264            // 348
        , -1.144    ,  0.088            // 349
        ,  -1.32    ,  0.264            // 350
        ,  -1.32    ,  0.088            // 351
        , -1.496    ,   1.32            // 352
        , -1.496    ,  1.144            // 353
        , -1.672    ,   1.32            // 354
        , -1.672    ,  1.144            // 355
        , -1.496    ,  0.968            // 356
        , -1.496    ,  0.792            // 357
        , -1.672    ,  0.968            // 358
        , -1.672    ,  0.792            // 359
        , -1.848    ,   1.32            // 360
        , -1.848    ,  1.144            // 361
        , -2.024    ,   1.32            // 362
        , -2.024    ,  1.144            // 363
        , -1.848    ,  0.968            // 364
        , -1.848    ,  0.792            // 365
        , -2.024    ,  0.968            // 366
        , -2.024    ,  0.792            // 367
        , -1.496    ,  0.616            // 368
        , -1.496    ,   0.44            // 369
        , -1.672    ,  0.616            // 370
        , -1.672    ,   0.44            // 371
        , -1.496    ,  0.264            // 372
        , -1.496    ,  0.088            // 373
        , -1.672    ,  0.264            // 374
        , -1.672    ,  0.088            // 375
        , -1.848    ,  0.616            // 376
        , -1.848    ,   0.44            // 377
        , -2.024    ,  0.616            // 378
        , -2.024    ,   0.44            // 379
        , -1.848    ,  0.264            // 380
        , -1.848    ,  0.088            // 381
        , -2.024    ,  0.264            // 382
        , -2.024    ,  0.088            // 383
        , -0.088    , -0.088            // 384
        , -0.088    , -0.264            // 385
        , -0.264    , -0.088            // 386
        , -0.264    , -0.264            // 387
        , -0.088    ,  -0.44            // 388
        , -0.088    , -0.616            // 389
        , -0.264    ,  -0.44            // 390
        , -0.264    , -0.616            // 391
        ,  -0.44    , -0.088            // 392
        ,  -0.44    , -0.264            // 393
        , -0.616    , -0.088            // 394
        , -0.616    , -0.264            // 395
        ,  -0.44    ,  -0.44            // 396
        ,  -0.44    , -0.616            // 397
        , -0.616    ,  -0.44            // 398
        , -0.616    , -0.616            // 399
        , -0.088    , -0.792            // 400
        , -0.088    , -0.968            // 401
        , -0.264    , -0.792            // 402
        , -0.264    , -0.968            // 403
        , -0.088    , -1.144            // 404
        , -0.088    ,  -1.32            // 405
        , -0.264    , -1.144            // 406
        , -0.264    ,  -1.32            // 407
        ,  -0.44    , -0.792            // 408
        ,  -0.44    , -0.968            // 409
        , -0.616    , -0.792            // 410
        , -0.616    , -0.968            // 411
        ,  -0.44    , -1.144            // 412
        ,  -0.44    ,  -1.32            // 413
        , -0.616    , -1.144            // 414
        , -0.616    ,  -1.32            // 415
        , -0.792    , -0.088            // 416
        , -0.792    , -0.264            // 417
        , -0.968    , -0.088            // 418
        , -0.968    , -0.264            // 419
        , -0.792    ,  -0.44            // 420
        , -0.792    , -0.616            // 421
        , -0.968    ,  -0.44            // 422
        , -0.968    , -0.616            // 423
        , -1.144    , -0.088            // 424
        , -1.144    , -0.264            // 425
        ,  -1.32    , -0.088            // 426
        ,  -1.32    , -0.264            // 427
        , -1.144    ,  -0.44            // 428
        , -1.144    , -0.616            // 429
        ,  -1.32    ,  -0.44            // 430
        ,  -1.32    , -0.616            // 431
        , -0.792    , -0.792            // 432
        , -0.792    , -0.968            // 433
        , -0.968    , -0.792            // 434
        , -0.968    , -0.968            // 435
        , -0.792    , -1.144            // 436
        , -0.792    ,  -1.32            // 437
        , -0.968    , -1.144            // 438
        , -0.968    ,  -1.32            // 439
        , -1.144    , -0.792            // 440
        , -1.144    , -0.968            // 441
        ,  -1.32    , -0.792            // 442
        ,  -1.32    , -0.968            // 443
        , -1.144    , -1.144            // 444
        , -1.144    ,  -1.32            // 445
        ,  -1.32    , -1.144            // 446
        ,  -1.32    ,  -1.32            // 447
        , -0.088    , -1.496            // 448
        , -0.088    , -1.672            // 449
        , -0.264    , -1.496            // 450
        , -0.264    , -1.672            // 451
        , -0.088    , -1.848            // 452
        , -0.088    , -2.024            // 453
        , -0.264    , -1.848            // 454
        , -0.264    , -2.024            // 455
        ,  -0.44    , -1.496            // 456
        ,  -0.44    , -1.672            // 457
        , -0.616    , -1.496            // 458
        , -0.616    , -1.672            // 459
        ,  -0.44    , -1.848            // 460
        ,  -0.44    , -2.024            // 461
        , -0.616    , -1.848            // 462
        , -0.616    , -2.024            // 463
        , -0.792    , -1.496            // 464
        , -0.792    , -1.672            // 465
        , -0.968    , -1.496            // 466
        , -0.968    , -1.672            // 467
        , -0.792    , -1.848            // 468
        , -0.792    , -2.024            // 469
        , -0.968    , -1.848            // 470
        , -0.968    , -2.024            // 471
        , -1.144    , -1.496            // 472
        , -1.144    , -1.672            // 473
        ,  -1.32    , -1.496            // 474
        ,  -1.32    , -1.672            // 475
        , -1.144    , -1.848            // 476
        , -1.144    , -2.024            // 477
        ,  -1.32    , -1.848            // 478
        ,  -1.32    , -2.024            // 479
        , -1.496    , -0.088            // 480
        , -1.496    , -0.264            // 481
        , -1.672    , -0.088            // 482
        , -1.672    , -0.264            // 483
        , -1.496    ,  -0.44            // 484
        , -1.496    , -0.616            // 485
        , -1.672    ,  -0.44            // 486
        , -1.672    , -0.616            // 487
        , -1.848    , -0.088            // 488
        , -1.848    , -0.264            // 489
        , -2.024    , -0.088            // 490
        , -2.024    , -0.264            // 491
        , -1.848    ,  -0.44            // 492
        , -1.848    , -0.616            // 493
        , -2.024    ,  -0.44            // 494
        , -2.024    , -0.616            // 495
        , -1.496    , -0.792            // 496
        , -1.496    , -0.968            // 497
        , -1.672    , -0.792            // 498
        , -1.672    , -0.968            // 499
        , -1.496    , -1.144            // 500
        , -1.496    ,  -1.32            // 501
        , -1.672    , -1.144            // 502
        , -1.672    ,  -1.32            // 503
        , -1.848    , -0.792            // 504
        , -1.848    , -0.968            // 505
        , -2.024    , -0.792            // 506
        , -2.024    , -0.968            // 507
        , -1.848    , -1.144            // 508
        , -1.848    ,  -1.32            // 509
        , -2.024    , -1.144            // 510
        , -2.024    ,  -1.32            // 511
    };