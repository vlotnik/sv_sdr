    DVBS2X_4_12_20_28APSK_132_180 : super.plane = {
            0.93    ,   0.93            // 0
        ,   0.93    ,  -0.93            // 1
        ,  -0.93    ,   0.93            // 2
        ,  -0.93    ,  -0.93            // 3
        ,  0.147    ,  1.306            // 4
        ,  0.147    , -1.306            // 5
        , -0.147    ,  1.306            // 6
        , -0.147    , -1.306            // 7
        ,  1.306    ,  0.147            // 8
        ,  1.306    , -0.147            // 9
        , -1.306    ,  0.147            // 10
        , -1.306    , -0.147            // 11
        ,  0.133    ,  0.133            // 12
        ,  0.133    , -0.133            // 13
        , -0.133    ,  0.133            // 14
        , -0.133    , -0.133            // 15
        ,  0.699    ,  1.113            // 16
        ,  0.699    , -1.113            // 17
        , -0.699    ,  1.113            // 18
        , -0.699    , -1.113            // 19
        ,  0.434    ,  1.241            // 20
        ,  0.434    , -1.241            // 21
        , -0.434    ,  1.241            // 22
        , -0.434    , -1.241            // 23
        ,  0.798    ,  0.126            // 24
        ,  0.798    , -0.126            // 25
        , -0.798    ,  0.126            // 26
        , -0.798    , -0.126            // 27
        ,  0.435    ,  0.117            // 28
        ,  0.435    , -0.117            // 29
        , -0.435    ,  0.117            // 30
        , -0.435    , -0.117            // 31
        ,  1.113    ,  0.699            // 32
        ,  1.113    , -0.699            // 33
        , -1.113    ,  0.699            // 34
        , -1.113    , -0.699            // 35
        ,  0.126    ,  0.798            // 36
        ,  0.126    , -0.798            // 37
        , -0.126    ,  0.798            // 38
        , -0.126    , -0.798            // 39
        ,  1.241    ,  0.434            // 40
        ,  1.241    , -0.434            // 41
        , -1.241    ,  0.434            // 42
        , -1.241    , -0.434            // 43
        ,  0.117    ,  0.435            // 44
        ,  0.117    , -0.435            // 45
        , -0.117    ,  0.435            // 46
        , -0.117    , -0.435            // 47
        ,  0.571    ,  0.571            // 48
        ,  0.571    , -0.571            // 49
        , -0.571    ,  0.571            // 50
        , -0.571    , -0.571            // 51
        ,  0.367    ,   0.72            // 52
        ,  0.367    ,  -0.72            // 53
        , -0.367    ,   0.72            // 54
        , -0.367    ,  -0.72            // 55
        ,   0.72    ,  0.367            // 56
        ,   0.72    , -0.367            // 57
        ,  -0.72    ,  0.367            // 58
        ,  -0.72    , -0.367            // 59
        ,  0.319    ,  0.319            // 60
        ,  0.319    , -0.319            // 61
        , -0.319    ,  0.319            // 62
        , -0.319    , -0.319            // 63
    };