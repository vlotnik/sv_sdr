    DVBS2X_256APSK_124_180 : super.plane = {
           0.259    ,  0.026            // 0
        ,  0.249    ,  0.076            // 1
        ,  0.201    ,  0.165            // 2
        ,   0.23    ,  0.123            // 3
        ,  0.026    ,  0.259            // 4
        ,  0.076    ,  0.249            // 5
        ,  0.165    ,  0.201            // 6
        ,  0.123    ,   0.23            // 7
        , -0.259    ,  0.026            // 8
        , -0.249    ,  0.076            // 9
        , -0.201    ,  0.165            // 10
        ,  -0.23    ,  0.123            // 11
        , -0.026    ,  0.259            // 12
        , -0.076    ,  0.249            // 13
        , -0.165    ,  0.201            // 14
        , -0.123    ,   0.23            // 15
        ,  0.259    , -0.026            // 16
        ,  0.249    , -0.076            // 17
        ,  0.201    , -0.165            // 18
        ,   0.23    , -0.123            // 19
        ,  0.026    , -0.259            // 20
        ,  0.076    , -0.249            // 21
        ,  0.165    , -0.201            // 22
        ,  0.123    ,  -0.23            // 23
        , -0.259    , -0.026            // 24
        , -0.249    , -0.076            // 25
        , -0.201    , -0.165            // 26
        ,  -0.23    , -0.123            // 27
        , -0.026    , -0.259            // 28
        , -0.076    , -0.249            // 29
        , -0.165    , -0.201            // 30
        , -0.123    ,  -0.23            // 31
        ,  0.464    ,  0.046            // 32
        ,  0.446    ,  0.135            // 33
        ,  0.361    ,  0.296            // 34
        ,  0.411    ,   0.22            // 35
        ,  0.046    ,  0.464            // 36
        ,  0.135    ,  0.446            // 37
        ,  0.296    ,  0.361            // 38
        ,   0.22    ,  0.411            // 39
        , -0.464    ,  0.046            // 40
        , -0.446    ,  0.135            // 41
        , -0.361    ,  0.296            // 42
        , -0.411    ,   0.22            // 43
        , -0.046    ,  0.464            // 44
        , -0.135    ,  0.446            // 45
        , -0.296    ,  0.361            // 46
        ,  -0.22    ,  0.411            // 47
        ,  0.464    , -0.046            // 48
        ,  0.446    , -0.135            // 49
        ,  0.361    , -0.296            // 50
        ,  0.411    ,  -0.22            // 51
        ,  0.046    , -0.464            // 52
        ,  0.135    , -0.446            // 53
        ,  0.296    , -0.361            // 54
        ,   0.22    , -0.411            // 55
        , -0.464    , -0.046            // 56
        , -0.446    , -0.135            // 57
        , -0.361    , -0.296            // 58
        , -0.411    ,  -0.22            // 59
        , -0.046    , -0.464            // 60
        , -0.135    , -0.446            // 61
        , -0.296    , -0.361            // 62
        ,  -0.22    , -0.411            // 63
        ,  0.772    ,  0.076            // 64
        ,  0.743    ,  0.225            // 65
        ,    0.6    ,  0.492            // 66
        ,  0.684    ,  0.366            // 67
        ,  0.076    ,  0.772            // 68
        ,  0.225    ,  0.743            // 69
        ,  0.492    ,    0.6            // 70
        ,  0.366    ,  0.684            // 71
        , -0.772    ,  0.076            // 72
        , -0.743    ,  0.225            // 73
        ,   -0.6    ,  0.492            // 74
        , -0.684    ,  0.366            // 75
        , -0.076    ,  0.772            // 76
        , -0.225    ,  0.743            // 77
        , -0.492    ,    0.6            // 78
        , -0.366    ,  0.684            // 79
        ,  0.772    , -0.076            // 80
        ,  0.743    , -0.225            // 81
        ,    0.6    , -0.492            // 82
        ,  0.684    , -0.366            // 83
        ,  0.076    , -0.772            // 84
        ,  0.225    , -0.743            // 85
        ,  0.492    ,   -0.6            // 86
        ,  0.366    , -0.684            // 87
        , -0.772    , -0.076            // 88
        , -0.743    , -0.225            // 89
        ,   -0.6    , -0.492            // 90
        , -0.684    , -0.366            // 91
        , -0.076    , -0.772            // 92
        , -0.225    , -0.743            // 93
        , -0.492    ,   -0.6            // 94
        , -0.366    , -0.684            // 95
        ,  0.623    ,  0.061            // 96
        ,  0.599    ,  0.182            // 97
        ,  0.484    ,  0.397            // 98
        ,  0.552    ,  0.295            // 99
        ,  0.061    ,  0.623            // 100
        ,  0.182    ,  0.599            // 101
        ,  0.397    ,  0.484            // 102
        ,  0.295    ,  0.552            // 103
        , -0.623    ,  0.061            // 104
        , -0.599    ,  0.182            // 105
        , -0.484    ,  0.397            // 106
        , -0.552    ,  0.295            // 107
        , -0.061    ,  0.623            // 108
        , -0.182    ,  0.599            // 109
        , -0.397    ,  0.484            // 110
        , -0.295    ,  0.552            // 111
        ,  0.623    , -0.061            // 112
        ,  0.599    , -0.182            // 113
        ,  0.484    , -0.397            // 114
        ,  0.552    , -0.295            // 115
        ,  0.061    , -0.623            // 116
        ,  0.182    , -0.599            // 117
        ,  0.397    , -0.484            // 118
        ,  0.295    , -0.552            // 119
        , -0.623    , -0.061            // 120
        , -0.599    , -0.182            // 121
        , -0.484    , -0.397            // 122
        , -0.552    , -0.295            // 123
        , -0.061    , -0.623            // 124
        , -0.182    , -0.599            // 125
        , -0.397    , -0.484            // 126
        , -0.295    , -0.552            // 127
        ,  1.694    ,  0.167            // 128
        ,  1.629    ,  0.494            // 129
        ,  1.316    ,   1.08            // 130
        ,  1.501    ,  0.802            // 131
        ,  0.167    ,  1.694            // 132
        ,  0.494    ,  1.629            // 133
        ,   1.08    ,  1.316            // 134
        ,  0.802    ,  1.501            // 135
        , -1.694    ,  0.167            // 136
        , -1.629    ,  0.494            // 137
        , -1.316    ,   1.08            // 138
        , -1.501    ,  0.802            // 139
        , -0.167    ,  1.694            // 140
        , -0.494    ,  1.629            // 141
        ,  -1.08    ,  1.316            // 142
        , -0.802    ,  1.501            // 143
        ,  1.694    , -0.167            // 144
        ,  1.629    , -0.494            // 145
        ,  1.316    ,  -1.08            // 146
        ,  1.501    , -0.802            // 147
        ,  0.167    , -1.694            // 148
        ,  0.494    , -1.629            // 149
        ,   1.08    , -1.316            // 150
        ,  0.802    , -1.501            // 151
        , -1.694    , -0.167            // 152
        , -1.629    , -0.494            // 153
        , -1.316    ,  -1.08            // 154
        , -1.501    , -0.802            // 155
        , -0.167    , -1.694            // 156
        , -0.494    , -1.629            // 157
        ,  -1.08    , -1.316            // 158
        , -0.802    , -1.501            // 159
        ,  1.316    ,   0.13            // 160
        ,  1.265    ,  0.384            // 161
        ,  1.022    ,  0.839            // 162
        ,  1.166    ,  0.623            // 163
        ,   0.13    ,  1.316            // 164
        ,  0.384    ,  1.265            // 165
        ,  0.839    ,  1.022            // 166
        ,  0.623    ,  1.166            // 167
        , -1.316    ,   0.13            // 168
        , -1.265    ,  0.384            // 169
        , -1.022    ,  0.839            // 170
        , -1.166    ,  0.623            // 171
        ,  -0.13    ,  1.316            // 172
        , -0.384    ,  1.265            // 173
        , -0.839    ,  1.022            // 174
        , -0.623    ,  1.166            // 175
        ,  1.316    ,  -0.13            // 176
        ,  1.265    , -0.384            // 177
        ,  1.022    , -0.839            // 178
        ,  1.166    , -0.623            // 179
        ,   0.13    , -1.316            // 180
        ,  0.384    , -1.265            // 181
        ,  0.839    , -1.022            // 182
        ,  0.623    , -1.166            // 183
        , -1.316    ,  -0.13            // 184
        , -1.265    , -0.384            // 185
        , -1.022    , -0.839            // 186
        , -1.166    , -0.623            // 187
        ,  -0.13    , -1.316            // 188
        , -0.384    , -1.265            // 189
        , -0.839    , -1.022            // 190
        , -0.623    , -1.166            // 191
        ,  0.925    ,  0.091            // 192
        ,  0.889    ,   0.27            // 193
        ,  0.718    ,   0.59            // 194
        ,   0.82    ,  0.438            // 195
        ,  0.091    ,  0.925            // 196
        ,   0.27    ,  0.889            // 197
        ,   0.59    ,  0.718            // 198
        ,  0.438    ,   0.82            // 199
        , -0.925    ,  0.091            // 200
        , -0.889    ,   0.27            // 201
        , -0.718    ,   0.59            // 202
        ,  -0.82    ,  0.438            // 203
        , -0.091    ,  0.925            // 204
        ,  -0.27    ,  0.889            // 205
        ,  -0.59    ,  0.718            // 206
        , -0.438    ,   0.82            // 207
        ,  0.925    , -0.091            // 208
        ,  0.889    ,  -0.27            // 209
        ,  0.718    ,  -0.59            // 210
        ,   0.82    , -0.438            // 211
        ,  0.091    , -0.925            // 212
        ,   0.27    , -0.889            // 213
        ,   0.59    , -0.718            // 214
        ,  0.438    ,  -0.82            // 215
        , -0.925    , -0.091            // 216
        , -0.889    ,  -0.27            // 217
        , -0.718    ,  -0.59            // 218
        ,  -0.82    , -0.438            // 219
        , -0.091    , -0.925            // 220
        ,  -0.27    , -0.889            // 221
        ,  -0.59    , -0.718            // 222
        , -0.438    ,  -0.82            // 223
        ,  1.097    ,  0.108            // 224
        ,  1.055    ,   0.32            // 225
        ,  0.852    ,    0.7            // 226
        ,  0.973    ,   0.52            // 227
        ,  0.108    ,  1.097            // 228
        ,   0.32    ,  1.055            // 229
        ,    0.7    ,  0.852            // 230
        ,   0.52    ,  0.973            // 231
        , -1.097    ,  0.108            // 232
        , -1.055    ,   0.32            // 233
        , -0.852    ,    0.7            // 234
        , -0.973    ,   0.52            // 235
        , -0.108    ,  1.097            // 236
        ,  -0.32    ,  1.055            // 237
        ,   -0.7    ,  0.852            // 238
        ,  -0.52    ,  0.973            // 239
        ,  1.097    , -0.108            // 240
        ,  1.055    ,  -0.32            // 241
        ,  0.852    ,   -0.7            // 242
        ,  0.973    ,  -0.52            // 243
        ,  0.108    , -1.097            // 244
        ,   0.32    , -1.055            // 245
        ,    0.7    , -0.852            // 246
        ,   0.52    , -0.973            // 247
        , -1.097    , -0.108            // 248
        , -1.055    ,  -0.32            // 249
        , -0.852    ,   -0.7            // 250
        , -0.973    ,  -0.52            // 251
        , -0.108    , -1.097            // 252
        ,  -0.32    , -1.055            // 253
        ,   -0.7    , -0.852            // 254
        ,  -0.52    , -0.973            // 255
    };