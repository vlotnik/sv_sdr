//--------------------------------------------------------------------------------------------------------------------------------
// name : raxi_bfm
//--------------------------------------------------------------------------------------------------------------------------------
interface raxi_bfm #(
      DW = pkg_raxi::RAXI_DEFAULT_DW
    , UW = pkg_raxi::RAXI_DEFAULT_UW
    , IW = pkg_raxi::RAXI_DEFAULT_IW
) (
      input clk
);
//--------------------------------------------------------------------------------------------------------------------------------
    bit                                 reset;
    bit                                 valid;
    bit                                 first;
    bit                                 last;
    bit                                 keep;
    bit                                 ready;
    bit[DW-1:0]                         data;
    bit[UW-1:0]                         user;
    bit[IW-1:0]                         id;
//--------------------------------------------------------------------------------------------------------------------------------
endinterface