    DVBS2X_4_12APSK_7_15 : super.plane = {
           0.804    ,  0.804            // 0
        ,  0.804    , -0.804            // 1
        , -0.804    ,  0.804            // 2
        , -0.804    , -0.804            // 3
        ,  1.099    ,  0.294            // 4
        ,  1.099    , -0.294            // 5
        , -1.099    ,  0.294            // 6
        , -1.099    , -0.294            // 7
        ,  0.294    ,  1.099            // 8
        ,  0.294    , -1.099            // 9
        , -0.294    ,  1.099            // 10
        , -0.294    , -1.099            // 11
        ,  0.242    ,  0.242            // 12
        ,  0.242    , -0.242            // 13
        , -0.242    ,  0.242            // 14
        , -0.242    , -0.242            // 15
    };