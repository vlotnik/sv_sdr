    DVBS2X_4_12APSK_28_45 : super.plane = {
           0.806    ,  0.806            // 0
        ,  0.806    , -0.806            // 1
        , -0.806    ,  0.806            // 2
        , -0.806    , -0.806            // 3
        ,    1.1    ,  0.295            // 4
        ,    1.1    , -0.295            // 5
        ,   -1.1    ,  0.295            // 6
        ,   -1.1    , -0.295            // 7
        ,  0.295    ,    1.1            // 8
        ,  0.295    ,   -1.1            // 9
        , -0.295    ,    1.1            // 10
        , -0.295    ,   -1.1            // 11
        ,   0.23    ,   0.23            // 12
        ,   0.23    ,  -0.23            // 13
        ,  -0.23    ,   0.23            // 14
        ,  -0.23    ,  -0.23            // 15
    };