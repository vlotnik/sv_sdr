    DVBS2X_8_8APSK_20_30 : super.plane = {
           0.506    ,  0.247            // 0
        ,  0.247    ,  0.506            // 1
        , -0.506    ,  0.247            // 2
        , -0.247    ,  0.506            // 3
        ,  0.506    , -0.247            // 4
        ,  0.247    , -0.506            // 5
        , -0.506    , -0.247            // 6
        , -0.247    , -0.506            // 7
        ,  1.201    ,  0.491            // 8
        ,  0.491    ,  1.201            // 9
        , -1.201    ,  0.491            // 10
        , -0.491    ,  1.201            // 11
        ,  1.201    , -0.491            // 12
        ,  0.491    , -1.201            // 13
        , -1.201    , -0.491            // 14
        , -0.491    , -1.201            // 15
    };