    DVBS2X_4_12_16RBAPSK_32_45 : super.plane = {
          -0.709    ,  1.061            // 0
        , -0.249    ,  1.252            // 1
        ,  0.709    ,  1.061            // 2
        ,  0.249    ,  1.252            // 3
        , -0.487    ,  0.487            // 4
        , -0.178    ,  0.666            // 5
        ,  0.487    ,  0.487            // 6
        ,  0.178    ,  0.666            // 7
        , -1.061    ,  0.709            // 8
        , -1.252    ,  0.249            // 9
        ,  1.061    ,  0.709            // 10
        ,  1.252    ,  0.249            // 11
        , -0.666    ,  0.178            // 12
        , -0.172    ,  0.172            // 13
        ,  0.666    ,  0.178            // 14
        ,  0.172    ,  0.172            // 15
        , -0.709    , -1.061            // 16
        , -0.249    , -1.252            // 17
        ,  0.709    , -1.061            // 18
        ,  0.249    , -1.252            // 19
        , -0.487    , -0.487            // 20
        , -0.178    , -0.666            // 21
        ,  0.487    , -0.487            // 22
        ,  0.178    , -0.666            // 23
        , -1.061    , -0.709            // 24
        , -1.252    , -0.249            // 25
        ,  1.061    , -0.709            // 26
        ,  1.252    , -0.249            // 27
        , -0.666    , -0.178            // 28
        , -0.172    , -0.172            // 29
        ,  0.666    , -0.178            // 30
        ,  0.172    , -0.172            // 31
    };