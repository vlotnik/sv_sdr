    DVBS2X_8_8APSK_96_180 : super.plane = {
           0.543    ,  0.225            // 0
        ,  0.225    ,  0.543            // 1
        , -0.543    ,  0.225            // 2
        , -0.225    ,  0.543            // 3
        ,  0.543    , -0.225            // 4
        ,  0.225    , -0.543            // 5
        , -0.543    , -0.225            // 6
        , -0.225    , -0.543            // 7
        ,  1.189    ,  0.492            // 8
        ,  0.492    ,  1.189            // 9
        , -1.189    ,  0.492            // 10
        , -0.492    ,  1.189            // 11
        ,  1.189    , -0.492            // 12
        ,  0.492    , -1.189            // 13
        , -1.189    , -0.492            // 14
        , -0.492    , -1.189            // 15
    };