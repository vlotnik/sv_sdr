    QAM128 : super.plane = {
           1.458    ,  0.928            // 0
        ,  1.458    ,  0.663            // 1
        ,  1.193    ,  0.928            // 2
        ,  1.193    ,  0.663            // 3
        ,  1.458    ,  0.398            // 4
        ,  1.458    ,  0.133            // 5
        ,  1.193    ,  0.398            // 6
        ,  1.193    ,  0.133            // 7
        ,  0.928    ,  1.458            // 8
        ,  0.928    ,  1.193            // 9
        ,  0.663    ,  1.458            // 10
        ,  0.663    ,  1.193            // 11
        ,  0.398    ,  1.458            // 12
        ,  0.398    ,  1.193            // 13
        ,  0.133    ,  1.458            // 14
        ,  0.133    ,  1.193            // 15
        ,  0.928    ,  0.928            // 16
        ,  0.928    ,  0.663            // 17
        ,  0.663    ,  0.928            // 18
        ,  0.663    ,  0.663            // 19
        ,  0.928    ,  0.398            // 20
        ,  0.928    ,  0.133            // 21
        ,  0.663    ,  0.398            // 22
        ,  0.663    ,  0.133            // 23
        ,  0.398    ,  0.928            // 24
        ,  0.398    ,  0.663            // 25
        ,  0.133    ,  0.928            // 26
        ,  0.133    ,  0.663            // 27
        ,  0.398    ,  0.398            // 28
        ,  0.398    ,  0.133            // 29
        ,  0.133    ,  0.398            // 30
        ,  0.133    ,  0.133            // 31
        ,  1.458    , -0.133            // 32
        ,  1.458    , -0.398            // 33
        ,  1.193    , -0.133            // 34
        ,  1.193    , -0.398            // 35
        ,  1.458    , -0.663            // 36
        ,  1.458    , -0.928            // 37
        ,  1.193    , -0.663            // 38
        ,  1.193    , -0.928            // 39
        ,  0.928    , -1.193            // 40
        ,  0.928    , -1.458            // 41
        ,  0.663    , -1.193            // 42
        ,  0.663    , -1.458            // 43
        ,  0.398    , -1.193            // 44
        ,  0.398    , -1.458            // 45
        ,  0.133    , -1.193            // 46
        ,  0.133    , -1.458            // 47
        ,  0.928    , -0.133            // 48
        ,  0.928    , -0.398            // 49
        ,  0.663    , -0.133            // 50
        ,  0.663    , -0.398            // 51
        ,  0.928    , -0.663            // 52
        ,  0.928    , -0.928            // 53
        ,  0.663    , -0.663            // 54
        ,  0.663    , -0.928            // 55
        ,  0.398    , -0.133            // 56
        ,  0.398    , -0.398            // 57
        ,  0.133    , -0.133            // 58
        ,  0.133    , -0.398            // 59
        ,  0.398    , -0.663            // 60
        ,  0.398    , -0.928            // 61
        ,  0.133    , -0.663            // 62
        ,  0.133    , -0.928            // 63
        , -0.133    ,  1.458            // 64
        , -0.133    ,  1.193            // 65
        , -0.398    ,  1.458            // 66
        , -0.398    ,  1.193            // 67
        , -0.663    ,  1.458            // 68
        , -0.663    ,  1.193            // 69
        , -0.928    ,  1.458            // 70
        , -0.928    ,  1.193            // 71
        , -1.193    ,  0.928            // 72
        , -1.193    ,  0.663            // 73
        , -1.458    ,  0.928            // 74
        , -1.458    ,  0.663            // 75
        , -1.193    ,  0.398            // 76
        , -1.193    ,  0.133            // 77
        , -1.458    ,  0.398            // 78
        , -1.458    ,  0.133            // 79
        , -0.133    ,  0.928            // 80
        , -0.133    ,  0.663            // 81
        , -0.398    ,  0.928            // 82
        , -0.398    ,  0.663            // 83
        , -0.133    ,  0.398            // 84
        , -0.133    ,  0.133            // 85
        , -0.398    ,  0.398            // 86
        , -0.398    ,  0.133            // 87
        , -0.663    ,  0.928            // 88
        , -0.663    ,  0.663            // 89
        , -0.928    ,  0.928            // 90
        , -0.928    ,  0.663            // 91
        , -0.663    ,  0.398            // 92
        , -0.663    ,  0.133            // 93
        , -0.928    ,  0.398            // 94
        , -0.928    ,  0.133            // 95
        , -0.133    , -1.193            // 96
        , -0.133    , -1.458            // 97
        , -0.398    , -1.193            // 98
        , -0.398    , -1.458            // 99
        , -0.663    , -1.193            // 100
        , -0.663    , -1.458            // 101
        , -0.928    , -1.193            // 102
        , -0.928    , -1.458            // 103
        , -1.193    , -0.133            // 104
        , -1.193    , -0.398            // 105
        , -1.458    , -0.133            // 106
        , -1.458    , -0.398            // 107
        , -1.193    , -0.663            // 108
        , -1.193    , -0.928            // 109
        , -1.458    , -0.663            // 110
        , -1.458    , -0.928            // 111
        , -0.133    , -0.133            // 112
        , -0.133    , -0.398            // 113
        , -0.398    , -0.133            // 114
        , -0.398    , -0.398            // 115
        , -0.133    , -0.663            // 116
        , -0.133    , -0.928            // 117
        , -0.398    , -0.663            // 118
        , -0.398    , -0.928            // 119
        , -0.663    , -0.133            // 120
        , -0.663    , -0.398            // 121
        , -0.928    , -0.133            // 122
        , -0.928    , -0.398            // 123
        , -0.663    , -0.663            // 124
        , -0.663    , -0.928            // 125
        , -0.928    , -0.663            // 126
        , -0.928    , -0.928            // 127
    };