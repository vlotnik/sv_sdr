    DVBS2X_4_12APSK_3_5 : super.plane = {
           0.807    ,  0.807            // 0
        ,  0.807    , -0.807            // 1
        , -0.807    ,  0.807            // 2
        , -0.807    , -0.807            // 3
        ,  1.102    ,  0.295            // 4
        ,  1.102    , -0.295            // 5
        , -1.102    ,  0.295            // 6
        , -1.102    , -0.295            // 7
        ,  0.295    ,  1.102            // 8
        ,  0.295    , -1.102            // 9
        , -0.295    ,  1.102            // 10
        , -0.295    , -1.102            // 11
        ,  0.218    ,  0.218            // 12
        ,  0.218    , -0.218            // 13
        , -0.218    ,  0.218            // 14
        , -0.218    , -0.218            // 15
    };