    QAM4096 : super.plane = {
           5.569    ,  5.569            // 0
        ,  5.569    ,  5.392            // 1
        ,  5.392    ,  5.569            // 2
        ,  5.392    ,  5.392            // 3
        ,  5.569    ,  5.039            // 4
        ,  5.569    ,  5.216            // 5
        ,  5.392    ,  5.039            // 6
        ,  5.392    ,  5.216            // 7
        ,  5.039    ,  5.569            // 8
        ,  5.039    ,  5.392            // 9
        ,  5.216    ,  5.569            // 10
        ,  5.216    ,  5.392            // 11
        ,  5.039    ,  5.039            // 12
        ,  5.039    ,  5.216            // 13
        ,  5.216    ,  5.039            // 14
        ,  5.216    ,  5.216            // 15
        ,  5.569    ,  4.332            // 16
        ,  5.569    ,  4.508            // 17
        ,  5.392    ,  4.332            // 18
        ,  5.392    ,  4.508            // 19
        ,  5.569    ,  4.862            // 20
        ,  5.569    ,  4.685            // 21
        ,  5.392    ,  4.862            // 22
        ,  5.392    ,  4.685            // 23
        ,  5.039    ,  4.332            // 24
        ,  5.039    ,  4.508            // 25
        ,  5.216    ,  4.332            // 26
        ,  5.216    ,  4.508            // 27
        ,  5.039    ,  4.862            // 28
        ,  5.039    ,  4.685            // 29
        ,  5.216    ,  4.862            // 30
        ,  5.216    ,  4.685            // 31
        ,  4.332    ,  5.569            // 32
        ,  4.332    ,  5.392            // 33
        ,  4.508    ,  5.569            // 34
        ,  4.508    ,  5.392            // 35
        ,  4.332    ,  5.039            // 36
        ,  4.332    ,  5.216            // 37
        ,  4.508    ,  5.039            // 38
        ,  4.508    ,  5.216            // 39
        ,  4.862    ,  5.569            // 40
        ,  4.862    ,  5.392            // 41
        ,  4.685    ,  5.569            // 42
        ,  4.685    ,  5.392            // 43
        ,  4.862    ,  5.039            // 44
        ,  4.862    ,  5.216            // 45
        ,  4.685    ,  5.039            // 46
        ,  4.685    ,  5.216            // 47
        ,  4.332    ,  4.332            // 48
        ,  4.332    ,  4.508            // 49
        ,  4.508    ,  4.332            // 50
        ,  4.508    ,  4.508            // 51
        ,  4.332    ,  4.862            // 52
        ,  4.332    ,  4.685            // 53
        ,  4.508    ,  4.862            // 54
        ,  4.508    ,  4.685            // 55
        ,  4.862    ,  4.332            // 56
        ,  4.862    ,  4.508            // 57
        ,  4.685    ,  4.332            // 58
        ,  4.685    ,  4.508            // 59
        ,  4.862    ,  4.862            // 60
        ,  4.862    ,  4.685            // 61
        ,  4.685    ,  4.862            // 62
        ,  4.685    ,  4.685            // 63
        ,  5.569    ,  2.917            // 64
        ,  5.569    ,  3.094            // 65
        ,  5.392    ,  2.917            // 66
        ,  5.392    ,  3.094            // 67
        ,  5.569    ,  3.448            // 68
        ,  5.569    ,  3.271            // 69
        ,  5.392    ,  3.448            // 70
        ,  5.392    ,  3.271            // 71
        ,  5.039    ,  2.917            // 72
        ,  5.039    ,  3.094            // 73
        ,  5.216    ,  2.917            // 74
        ,  5.216    ,  3.094            // 75
        ,  5.039    ,  3.448            // 76
        ,  5.039    ,  3.271            // 77
        ,  5.216    ,  3.448            // 78
        ,  5.216    ,  3.271            // 79
        ,  5.569    ,  4.155            // 80
        ,  5.569    ,  3.978            // 81
        ,  5.392    ,  4.155            // 82
        ,  5.392    ,  3.978            // 83
        ,  5.569    ,  3.624            // 84
        ,  5.569    ,  3.801            // 85
        ,  5.392    ,  3.624            // 86
        ,  5.392    ,  3.801            // 87
        ,  5.039    ,  4.155            // 88
        ,  5.039    ,  3.978            // 89
        ,  5.216    ,  4.155            // 90
        ,  5.216    ,  3.978            // 91
        ,  5.039    ,  3.624            // 92
        ,  5.039    ,  3.801            // 93
        ,  5.216    ,  3.624            // 94
        ,  5.216    ,  3.801            // 95
        ,  4.332    ,  2.917            // 96
        ,  4.332    ,  3.094            // 97
        ,  4.508    ,  2.917            // 98
        ,  4.508    ,  3.094            // 99
        ,  4.332    ,  3.448            // 100
        ,  4.332    ,  3.271            // 101
        ,  4.508    ,  3.448            // 102
        ,  4.508    ,  3.271            // 103
        ,  4.862    ,  2.917            // 104
        ,  4.862    ,  3.094            // 105
        ,  4.685    ,  2.917            // 106
        ,  4.685    ,  3.094            // 107
        ,  4.862    ,  3.448            // 108
        ,  4.862    ,  3.271            // 109
        ,  4.685    ,  3.448            // 110
        ,  4.685    ,  3.271            // 111
        ,  4.332    ,  4.155            // 112
        ,  4.332    ,  3.978            // 113
        ,  4.508    ,  4.155            // 114
        ,  4.508    ,  3.978            // 115
        ,  4.332    ,  3.624            // 116
        ,  4.332    ,  3.801            // 117
        ,  4.508    ,  3.624            // 118
        ,  4.508    ,  3.801            // 119
        ,  4.862    ,  4.155            // 120
        ,  4.862    ,  3.978            // 121
        ,  4.685    ,  4.155            // 122
        ,  4.685    ,  3.978            // 123
        ,  4.862    ,  3.624            // 124
        ,  4.862    ,  3.801            // 125
        ,  4.685    ,  3.624            // 126
        ,  4.685    ,  3.801            // 127
        ,  2.917    ,  5.569            // 128
        ,  2.917    ,  5.392            // 129
        ,  3.094    ,  5.569            // 130
        ,  3.094    ,  5.392            // 131
        ,  2.917    ,  5.039            // 132
        ,  2.917    ,  5.216            // 133
        ,  3.094    ,  5.039            // 134
        ,  3.094    ,  5.216            // 135
        ,  3.448    ,  5.569            // 136
        ,  3.448    ,  5.392            // 137
        ,  3.271    ,  5.569            // 138
        ,  3.271    ,  5.392            // 139
        ,  3.448    ,  5.039            // 140
        ,  3.448    ,  5.216            // 141
        ,  3.271    ,  5.039            // 142
        ,  3.271    ,  5.216            // 143
        ,  2.917    ,  4.332            // 144
        ,  2.917    ,  4.508            // 145
        ,  3.094    ,  4.332            // 146
        ,  3.094    ,  4.508            // 147
        ,  2.917    ,  4.862            // 148
        ,  2.917    ,  4.685            // 149
        ,  3.094    ,  4.862            // 150
        ,  3.094    ,  4.685            // 151
        ,  3.448    ,  4.332            // 152
        ,  3.448    ,  4.508            // 153
        ,  3.271    ,  4.332            // 154
        ,  3.271    ,  4.508            // 155
        ,  3.448    ,  4.862            // 156
        ,  3.448    ,  4.685            // 157
        ,  3.271    ,  4.862            // 158
        ,  3.271    ,  4.685            // 159
        ,  4.155    ,  5.569            // 160
        ,  4.155    ,  5.392            // 161
        ,  3.978    ,  5.569            // 162
        ,  3.978    ,  5.392            // 163
        ,  4.155    ,  5.039            // 164
        ,  4.155    ,  5.216            // 165
        ,  3.978    ,  5.039            // 166
        ,  3.978    ,  5.216            // 167
        ,  3.624    ,  5.569            // 168
        ,  3.624    ,  5.392            // 169
        ,  3.801    ,  5.569            // 170
        ,  3.801    ,  5.392            // 171
        ,  3.624    ,  5.039            // 172
        ,  3.624    ,  5.216            // 173
        ,  3.801    ,  5.039            // 174
        ,  3.801    ,  5.216            // 175
        ,  4.155    ,  4.332            // 176
        ,  4.155    ,  4.508            // 177
        ,  3.978    ,  4.332            // 178
        ,  3.978    ,  4.508            // 179
        ,  4.155    ,  4.862            // 180
        ,  4.155    ,  4.685            // 181
        ,  3.978    ,  4.862            // 182
        ,  3.978    ,  4.685            // 183
        ,  3.624    ,  4.332            // 184
        ,  3.624    ,  4.508            // 185
        ,  3.801    ,  4.332            // 186
        ,  3.801    ,  4.508            // 187
        ,  3.624    ,  4.862            // 188
        ,  3.624    ,  4.685            // 189
        ,  3.801    ,  4.862            // 190
        ,  3.801    ,  4.685            // 191
        ,  2.917    ,  2.917            // 192
        ,  2.917    ,  3.094            // 193
        ,  3.094    ,  2.917            // 194
        ,  3.094    ,  3.094            // 195
        ,  2.917    ,  3.448            // 196
        ,  2.917    ,  3.271            // 197
        ,  3.094    ,  3.448            // 198
        ,  3.094    ,  3.271            // 199
        ,  3.448    ,  2.917            // 200
        ,  3.448    ,  3.094            // 201
        ,  3.271    ,  2.917            // 202
        ,  3.271    ,  3.094            // 203
        ,  3.448    ,  3.448            // 204
        ,  3.448    ,  3.271            // 205
        ,  3.271    ,  3.448            // 206
        ,  3.271    ,  3.271            // 207
        ,  2.917    ,  4.155            // 208
        ,  2.917    ,  3.978            // 209
        ,  3.094    ,  4.155            // 210
        ,  3.094    ,  3.978            // 211
        ,  2.917    ,  3.624            // 212
        ,  2.917    ,  3.801            // 213
        ,  3.094    ,  3.624            // 214
        ,  3.094    ,  3.801            // 215
        ,  3.448    ,  4.155            // 216
        ,  3.448    ,  3.978            // 217
        ,  3.271    ,  4.155            // 218
        ,  3.271    ,  3.978            // 219
        ,  3.448    ,  3.624            // 220
        ,  3.448    ,  3.801            // 221
        ,  3.271    ,  3.624            // 222
        ,  3.271    ,  3.801            // 223
        ,  4.155    ,  2.917            // 224
        ,  4.155    ,  3.094            // 225
        ,  3.978    ,  2.917            // 226
        ,  3.978    ,  3.094            // 227
        ,  4.155    ,  3.448            // 228
        ,  4.155    ,  3.271            // 229
        ,  3.978    ,  3.448            // 230
        ,  3.978    ,  3.271            // 231
        ,  3.624    ,  2.917            // 232
        ,  3.624    ,  3.094            // 233
        ,  3.801    ,  2.917            // 234
        ,  3.801    ,  3.094            // 235
        ,  3.624    ,  3.448            // 236
        ,  3.624    ,  3.271            // 237
        ,  3.801    ,  3.448            // 238
        ,  3.801    ,  3.271            // 239
        ,  4.155    ,  4.155            // 240
        ,  4.155    ,  3.978            // 241
        ,  3.978    ,  4.155            // 242
        ,  3.978    ,  3.978            // 243
        ,  4.155    ,  3.624            // 244
        ,  4.155    ,  3.801            // 245
        ,  3.978    ,  3.624            // 246
        ,  3.978    ,  3.801            // 247
        ,  3.624    ,  4.155            // 248
        ,  3.624    ,  3.978            // 249
        ,  3.801    ,  4.155            // 250
        ,  3.801    ,  3.978            // 251
        ,  3.624    ,  3.624            // 252
        ,  3.624    ,  3.801            // 253
        ,  3.801    ,  3.624            // 254
        ,  3.801    ,  3.801            // 255
        ,  5.569    ,  0.088            // 256
        ,  5.569    ,  0.265            // 257
        ,  5.392    ,  0.088            // 258
        ,  5.392    ,  0.265            // 259
        ,  5.569    ,  0.619            // 260
        ,  5.569    ,  0.442            // 261
        ,  5.392    ,  0.619            // 262
        ,  5.392    ,  0.442            // 263
        ,  5.039    ,  0.088            // 264
        ,  5.039    ,  0.265            // 265
        ,  5.216    ,  0.088            // 266
        ,  5.216    ,  0.265            // 267
        ,  5.039    ,  0.619            // 268
        ,  5.039    ,  0.442            // 269
        ,  5.216    ,  0.619            // 270
        ,  5.216    ,  0.442            // 271
        ,  5.569    ,  1.326            // 272
        ,  5.569    ,  1.149            // 273
        ,  5.392    ,  1.326            // 274
        ,  5.392    ,  1.149            // 275
        ,  5.569    ,  0.796            // 276
        ,  5.569    ,  0.972            // 277
        ,  5.392    ,  0.796            // 278
        ,  5.392    ,  0.972            // 279
        ,  5.039    ,  1.326            // 280
        ,  5.039    ,  1.149            // 281
        ,  5.216    ,  1.326            // 282
        ,  5.216    ,  1.149            // 283
        ,  5.039    ,  0.796            // 284
        ,  5.039    ,  0.972            // 285
        ,  5.216    ,  0.796            // 286
        ,  5.216    ,  0.972            // 287
        ,  4.332    ,  0.088            // 288
        ,  4.332    ,  0.265            // 289
        ,  4.508    ,  0.088            // 290
        ,  4.508    ,  0.265            // 291
        ,  4.332    ,  0.619            // 292
        ,  4.332    ,  0.442            // 293
        ,  4.508    ,  0.619            // 294
        ,  4.508    ,  0.442            // 295
        ,  4.862    ,  0.088            // 296
        ,  4.862    ,  0.265            // 297
        ,  4.685    ,  0.088            // 298
        ,  4.685    ,  0.265            // 299
        ,  4.862    ,  0.619            // 300
        ,  4.862    ,  0.442            // 301
        ,  4.685    ,  0.619            // 302
        ,  4.685    ,  0.442            // 303
        ,  4.332    ,  1.326            // 304
        ,  4.332    ,  1.149            // 305
        ,  4.508    ,  1.326            // 306
        ,  4.508    ,  1.149            // 307
        ,  4.332    ,  0.796            // 308
        ,  4.332    ,  0.972            // 309
        ,  4.508    ,  0.796            // 310
        ,  4.508    ,  0.972            // 311
        ,  4.862    ,  1.326            // 312
        ,  4.862    ,  1.149            // 313
        ,  4.685    ,  1.326            // 314
        ,  4.685    ,  1.149            // 315
        ,  4.862    ,  0.796            // 316
        ,  4.862    ,  0.972            // 317
        ,  4.685    ,  0.796            // 318
        ,  4.685    ,  0.972            // 319
        ,  5.569    ,   2.74            // 320
        ,  5.569    ,  2.564            // 321
        ,  5.392    ,   2.74            // 322
        ,  5.392    ,  2.564            // 323
        ,  5.569    ,   2.21            // 324
        ,  5.569    ,  2.387            // 325
        ,  5.392    ,   2.21            // 326
        ,  5.392    ,  2.387            // 327
        ,  5.039    ,   2.74            // 328
        ,  5.039    ,  2.564            // 329
        ,  5.216    ,   2.74            // 330
        ,  5.216    ,  2.564            // 331
        ,  5.039    ,   2.21            // 332
        ,  5.039    ,  2.387            // 333
        ,  5.216    ,   2.21            // 334
        ,  5.216    ,  2.387            // 335
        ,  5.569    ,  1.503            // 336
        ,  5.569    ,   1.68            // 337
        ,  5.392    ,  1.503            // 338
        ,  5.392    ,   1.68            // 339
        ,  5.569    ,  2.033            // 340
        ,  5.569    ,  1.856            // 341
        ,  5.392    ,  2.033            // 342
        ,  5.392    ,  1.856            // 343
        ,  5.039    ,  1.503            // 344
        ,  5.039    ,   1.68            // 345
        ,  5.216    ,  1.503            // 346
        ,  5.216    ,   1.68            // 347
        ,  5.039    ,  2.033            // 348
        ,  5.039    ,  1.856            // 349
        ,  5.216    ,  2.033            // 350
        ,  5.216    ,  1.856            // 351
        ,  4.332    ,   2.74            // 352
        ,  4.332    ,  2.564            // 353
        ,  4.508    ,   2.74            // 354
        ,  4.508    ,  2.564            // 355
        ,  4.332    ,   2.21            // 356
        ,  4.332    ,  2.387            // 357
        ,  4.508    ,   2.21            // 358
        ,  4.508    ,  2.387            // 359
        ,  4.862    ,   2.74            // 360
        ,  4.862    ,  2.564            // 361
        ,  4.685    ,   2.74            // 362
        ,  4.685    ,  2.564            // 363
        ,  4.862    ,   2.21            // 364
        ,  4.862    ,  2.387            // 365
        ,  4.685    ,   2.21            // 366
        ,  4.685    ,  2.387            // 367
        ,  4.332    ,  1.503            // 368
        ,  4.332    ,   1.68            // 369
        ,  4.508    ,  1.503            // 370
        ,  4.508    ,   1.68            // 371
        ,  4.332    ,  2.033            // 372
        ,  4.332    ,  1.856            // 373
        ,  4.508    ,  2.033            // 374
        ,  4.508    ,  1.856            // 375
        ,  4.862    ,  1.503            // 376
        ,  4.862    ,   1.68            // 377
        ,  4.685    ,  1.503            // 378
        ,  4.685    ,   1.68            // 379
        ,  4.862    ,  2.033            // 380
        ,  4.862    ,  1.856            // 381
        ,  4.685    ,  2.033            // 382
        ,  4.685    ,  1.856            // 383
        ,  2.917    ,  0.088            // 384
        ,  2.917    ,  0.265            // 385
        ,  3.094    ,  0.088            // 386
        ,  3.094    ,  0.265            // 387
        ,  2.917    ,  0.619            // 388
        ,  2.917    ,  0.442            // 389
        ,  3.094    ,  0.619            // 390
        ,  3.094    ,  0.442            // 391
        ,  3.448    ,  0.088            // 392
        ,  3.448    ,  0.265            // 393
        ,  3.271    ,  0.088            // 394
        ,  3.271    ,  0.265            // 395
        ,  3.448    ,  0.619            // 396
        ,  3.448    ,  0.442            // 397
        ,  3.271    ,  0.619            // 398
        ,  3.271    ,  0.442            // 399
        ,  2.917    ,  1.326            // 400
        ,  2.917    ,  1.149            // 401
        ,  3.094    ,  1.326            // 402
        ,  3.094    ,  1.149            // 403
        ,  2.917    ,  0.796            // 404
        ,  2.917    ,  0.972            // 405
        ,  3.094    ,  0.796            // 406
        ,  3.094    ,  0.972            // 407
        ,  3.448    ,  1.326            // 408
        ,  3.448    ,  1.149            // 409
        ,  3.271    ,  1.326            // 410
        ,  3.271    ,  1.149            // 411
        ,  3.448    ,  0.796            // 412
        ,  3.448    ,  0.972            // 413
        ,  3.271    ,  0.796            // 414
        ,  3.271    ,  0.972            // 415
        ,  4.155    ,  0.088            // 416
        ,  4.155    ,  0.265            // 417
        ,  3.978    ,  0.088            // 418
        ,  3.978    ,  0.265            // 419
        ,  4.155    ,  0.619            // 420
        ,  4.155    ,  0.442            // 421
        ,  3.978    ,  0.619            // 422
        ,  3.978    ,  0.442            // 423
        ,  3.624    ,  0.088            // 424
        ,  3.624    ,  0.265            // 425
        ,  3.801    ,  0.088            // 426
        ,  3.801    ,  0.265            // 427
        ,  3.624    ,  0.619            // 428
        ,  3.624    ,  0.442            // 429
        ,  3.801    ,  0.619            // 430
        ,  3.801    ,  0.442            // 431
        ,  4.155    ,  1.326            // 432
        ,  4.155    ,  1.149            // 433
        ,  3.978    ,  1.326            // 434
        ,  3.978    ,  1.149            // 435
        ,  4.155    ,  0.796            // 436
        ,  4.155    ,  0.972            // 437
        ,  3.978    ,  0.796            // 438
        ,  3.978    ,  0.972            // 439
        ,  3.624    ,  1.326            // 440
        ,  3.624    ,  1.149            // 441
        ,  3.801    ,  1.326            // 442
        ,  3.801    ,  1.149            // 443
        ,  3.624    ,  0.796            // 444
        ,  3.624    ,  0.972            // 445
        ,  3.801    ,  0.796            // 446
        ,  3.801    ,  0.972            // 447
        ,  2.917    ,   2.74            // 448
        ,  2.917    ,  2.564            // 449
        ,  3.094    ,   2.74            // 450
        ,  3.094    ,  2.564            // 451
        ,  2.917    ,   2.21            // 452
        ,  2.917    ,  2.387            // 453
        ,  3.094    ,   2.21            // 454
        ,  3.094    ,  2.387            // 455
        ,  3.448    ,   2.74            // 456
        ,  3.448    ,  2.564            // 457
        ,  3.271    ,   2.74            // 458
        ,  3.271    ,  2.564            // 459
        ,  3.448    ,   2.21            // 460
        ,  3.448    ,  2.387            // 461
        ,  3.271    ,   2.21            // 462
        ,  3.271    ,  2.387            // 463
        ,  2.917    ,  1.503            // 464
        ,  2.917    ,   1.68            // 465
        ,  3.094    ,  1.503            // 466
        ,  3.094    ,   1.68            // 467
        ,  2.917    ,  2.033            // 468
        ,  2.917    ,  1.856            // 469
        ,  3.094    ,  2.033            // 470
        ,  3.094    ,  1.856            // 471
        ,  3.448    ,  1.503            // 472
        ,  3.448    ,   1.68            // 473
        ,  3.271    ,  1.503            // 474
        ,  3.271    ,   1.68            // 475
        ,  3.448    ,  2.033            // 476
        ,  3.448    ,  1.856            // 477
        ,  3.271    ,  2.033            // 478
        ,  3.271    ,  1.856            // 479
        ,  4.155    ,   2.74            // 480
        ,  4.155    ,  2.564            // 481
        ,  3.978    ,   2.74            // 482
        ,  3.978    ,  2.564            // 483
        ,  4.155    ,   2.21            // 484
        ,  4.155    ,  2.387            // 485
        ,  3.978    ,   2.21            // 486
        ,  3.978    ,  2.387            // 487
        ,  3.624    ,   2.74            // 488
        ,  3.624    ,  2.564            // 489
        ,  3.801    ,   2.74            // 490
        ,  3.801    ,  2.564            // 491
        ,  3.624    ,   2.21            // 492
        ,  3.624    ,  2.387            // 493
        ,  3.801    ,   2.21            // 494
        ,  3.801    ,  2.387            // 495
        ,  4.155    ,  1.503            // 496
        ,  4.155    ,   1.68            // 497
        ,  3.978    ,  1.503            // 498
        ,  3.978    ,   1.68            // 499
        ,  4.155    ,  2.033            // 500
        ,  4.155    ,  1.856            // 501
        ,  3.978    ,  2.033            // 502
        ,  3.978    ,  1.856            // 503
        ,  3.624    ,  1.503            // 504
        ,  3.624    ,   1.68            // 505
        ,  3.801    ,  1.503            // 506
        ,  3.801    ,   1.68            // 507
        ,  3.624    ,  2.033            // 508
        ,  3.624    ,  1.856            // 509
        ,  3.801    ,  2.033            // 510
        ,  3.801    ,  1.856            // 511
        ,  0.088    ,  5.569            // 512
        ,  0.088    ,  5.392            // 513
        ,  0.265    ,  5.569            // 514
        ,  0.265    ,  5.392            // 515
        ,  0.088    ,  5.039            // 516
        ,  0.088    ,  5.216            // 517
        ,  0.265    ,  5.039            // 518
        ,  0.265    ,  5.216            // 519
        ,  0.619    ,  5.569            // 520
        ,  0.619    ,  5.392            // 521
        ,  0.442    ,  5.569            // 522
        ,  0.442    ,  5.392            // 523
        ,  0.619    ,  5.039            // 524
        ,  0.619    ,  5.216            // 525
        ,  0.442    ,  5.039            // 526
        ,  0.442    ,  5.216            // 527
        ,  0.088    ,  4.332            // 528
        ,  0.088    ,  4.508            // 529
        ,  0.265    ,  4.332            // 530
        ,  0.265    ,  4.508            // 531
        ,  0.088    ,  4.862            // 532
        ,  0.088    ,  4.685            // 533
        ,  0.265    ,  4.862            // 534
        ,  0.265    ,  4.685            // 535
        ,  0.619    ,  4.332            // 536
        ,  0.619    ,  4.508            // 537
        ,  0.442    ,  4.332            // 538
        ,  0.442    ,  4.508            // 539
        ,  0.619    ,  4.862            // 540
        ,  0.619    ,  4.685            // 541
        ,  0.442    ,  4.862            // 542
        ,  0.442    ,  4.685            // 543
        ,  1.326    ,  5.569            // 544
        ,  1.326    ,  5.392            // 545
        ,  1.149    ,  5.569            // 546
        ,  1.149    ,  5.392            // 547
        ,  1.326    ,  5.039            // 548
        ,  1.326    ,  5.216            // 549
        ,  1.149    ,  5.039            // 550
        ,  1.149    ,  5.216            // 551
        ,  0.796    ,  5.569            // 552
        ,  0.796    ,  5.392            // 553
        ,  0.972    ,  5.569            // 554
        ,  0.972    ,  5.392            // 555
        ,  0.796    ,  5.039            // 556
        ,  0.796    ,  5.216            // 557
        ,  0.972    ,  5.039            // 558
        ,  0.972    ,  5.216            // 559
        ,  1.326    ,  4.332            // 560
        ,  1.326    ,  4.508            // 561
        ,  1.149    ,  4.332            // 562
        ,  1.149    ,  4.508            // 563
        ,  1.326    ,  4.862            // 564
        ,  1.326    ,  4.685            // 565
        ,  1.149    ,  4.862            // 566
        ,  1.149    ,  4.685            // 567
        ,  0.796    ,  4.332            // 568
        ,  0.796    ,  4.508            // 569
        ,  0.972    ,  4.332            // 570
        ,  0.972    ,  4.508            // 571
        ,  0.796    ,  4.862            // 572
        ,  0.796    ,  4.685            // 573
        ,  0.972    ,  4.862            // 574
        ,  0.972    ,  4.685            // 575
        ,  0.088    ,  2.917            // 576
        ,  0.088    ,  3.094            // 577
        ,  0.265    ,  2.917            // 578
        ,  0.265    ,  3.094            // 579
        ,  0.088    ,  3.448            // 580
        ,  0.088    ,  3.271            // 581
        ,  0.265    ,  3.448            // 582
        ,  0.265    ,  3.271            // 583
        ,  0.619    ,  2.917            // 584
        ,  0.619    ,  3.094            // 585
        ,  0.442    ,  2.917            // 586
        ,  0.442    ,  3.094            // 587
        ,  0.619    ,  3.448            // 588
        ,  0.619    ,  3.271            // 589
        ,  0.442    ,  3.448            // 590
        ,  0.442    ,  3.271            // 591
        ,  0.088    ,  4.155            // 592
        ,  0.088    ,  3.978            // 593
        ,  0.265    ,  4.155            // 594
        ,  0.265    ,  3.978            // 595
        ,  0.088    ,  3.624            // 596
        ,  0.088    ,  3.801            // 597
        ,  0.265    ,  3.624            // 598
        ,  0.265    ,  3.801            // 599
        ,  0.619    ,  4.155            // 600
        ,  0.619    ,  3.978            // 601
        ,  0.442    ,  4.155            // 602
        ,  0.442    ,  3.978            // 603
        ,  0.619    ,  3.624            // 604
        ,  0.619    ,  3.801            // 605
        ,  0.442    ,  3.624            // 606
        ,  0.442    ,  3.801            // 607
        ,  1.326    ,  2.917            // 608
        ,  1.326    ,  3.094            // 609
        ,  1.149    ,  2.917            // 610
        ,  1.149    ,  3.094            // 611
        ,  1.326    ,  3.448            // 612
        ,  1.326    ,  3.271            // 613
        ,  1.149    ,  3.448            // 614
        ,  1.149    ,  3.271            // 615
        ,  0.796    ,  2.917            // 616
        ,  0.796    ,  3.094            // 617
        ,  0.972    ,  2.917            // 618
        ,  0.972    ,  3.094            // 619
        ,  0.796    ,  3.448            // 620
        ,  0.796    ,  3.271            // 621
        ,  0.972    ,  3.448            // 622
        ,  0.972    ,  3.271            // 623
        ,  1.326    ,  4.155            // 624
        ,  1.326    ,  3.978            // 625
        ,  1.149    ,  4.155            // 626
        ,  1.149    ,  3.978            // 627
        ,  1.326    ,  3.624            // 628
        ,  1.326    ,  3.801            // 629
        ,  1.149    ,  3.624            // 630
        ,  1.149    ,  3.801            // 631
        ,  0.796    ,  4.155            // 632
        ,  0.796    ,  3.978            // 633
        ,  0.972    ,  4.155            // 634
        ,  0.972    ,  3.978            // 635
        ,  0.796    ,  3.624            // 636
        ,  0.796    ,  3.801            // 637
        ,  0.972    ,  3.624            // 638
        ,  0.972    ,  3.801            // 639
        ,   2.74    ,  5.569            // 640
        ,   2.74    ,  5.392            // 641
        ,  2.564    ,  5.569            // 642
        ,  2.564    ,  5.392            // 643
        ,   2.74    ,  5.039            // 644
        ,   2.74    ,  5.216            // 645
        ,  2.564    ,  5.039            // 646
        ,  2.564    ,  5.216            // 647
        ,   2.21    ,  5.569            // 648
        ,   2.21    ,  5.392            // 649
        ,  2.387    ,  5.569            // 650
        ,  2.387    ,  5.392            // 651
        ,   2.21    ,  5.039            // 652
        ,   2.21    ,  5.216            // 653
        ,  2.387    ,  5.039            // 654
        ,  2.387    ,  5.216            // 655
        ,   2.74    ,  4.332            // 656
        ,   2.74    ,  4.508            // 657
        ,  2.564    ,  4.332            // 658
        ,  2.564    ,  4.508            // 659
        ,   2.74    ,  4.862            // 660
        ,   2.74    ,  4.685            // 661
        ,  2.564    ,  4.862            // 662
        ,  2.564    ,  4.685            // 663
        ,   2.21    ,  4.332            // 664
        ,   2.21    ,  4.508            // 665
        ,  2.387    ,  4.332            // 666
        ,  2.387    ,  4.508            // 667
        ,   2.21    ,  4.862            // 668
        ,   2.21    ,  4.685            // 669
        ,  2.387    ,  4.862            // 670
        ,  2.387    ,  4.685            // 671
        ,  1.503    ,  5.569            // 672
        ,  1.503    ,  5.392            // 673
        ,   1.68    ,  5.569            // 674
        ,   1.68    ,  5.392            // 675
        ,  1.503    ,  5.039            // 676
        ,  1.503    ,  5.216            // 677
        ,   1.68    ,  5.039            // 678
        ,   1.68    ,  5.216            // 679
        ,  2.033    ,  5.569            // 680
        ,  2.033    ,  5.392            // 681
        ,  1.856    ,  5.569            // 682
        ,  1.856    ,  5.392            // 683
        ,  2.033    ,  5.039            // 684
        ,  2.033    ,  5.216            // 685
        ,  1.856    ,  5.039            // 686
        ,  1.856    ,  5.216            // 687
        ,  1.503    ,  4.332            // 688
        ,  1.503    ,  4.508            // 689
        ,   1.68    ,  4.332            // 690
        ,   1.68    ,  4.508            // 691
        ,  1.503    ,  4.862            // 692
        ,  1.503    ,  4.685            // 693
        ,   1.68    ,  4.862            // 694
        ,   1.68    ,  4.685            // 695
        ,  2.033    ,  4.332            // 696
        ,  2.033    ,  4.508            // 697
        ,  1.856    ,  4.332            // 698
        ,  1.856    ,  4.508            // 699
        ,  2.033    ,  4.862            // 700
        ,  2.033    ,  4.685            // 701
        ,  1.856    ,  4.862            // 702
        ,  1.856    ,  4.685            // 703
        ,   2.74    ,  2.917            // 704
        ,   2.74    ,  3.094            // 705
        ,  2.564    ,  2.917            // 706
        ,  2.564    ,  3.094            // 707
        ,   2.74    ,  3.448            // 708
        ,   2.74    ,  3.271            // 709
        ,  2.564    ,  3.448            // 710
        ,  2.564    ,  3.271            // 711
        ,   2.21    ,  2.917            // 712
        ,   2.21    ,  3.094            // 713
        ,  2.387    ,  2.917            // 714
        ,  2.387    ,  3.094            // 715
        ,   2.21    ,  3.448            // 716
        ,   2.21    ,  3.271            // 717
        ,  2.387    ,  3.448            // 718
        ,  2.387    ,  3.271            // 719
        ,   2.74    ,  4.155            // 720
        ,   2.74    ,  3.978            // 721
        ,  2.564    ,  4.155            // 722
        ,  2.564    ,  3.978            // 723
        ,   2.74    ,  3.624            // 724
        ,   2.74    ,  3.801            // 725
        ,  2.564    ,  3.624            // 726
        ,  2.564    ,  3.801            // 727
        ,   2.21    ,  4.155            // 728
        ,   2.21    ,  3.978            // 729
        ,  2.387    ,  4.155            // 730
        ,  2.387    ,  3.978            // 731
        ,   2.21    ,  3.624            // 732
        ,   2.21    ,  3.801            // 733
        ,  2.387    ,  3.624            // 734
        ,  2.387    ,  3.801            // 735
        ,  1.503    ,  2.917            // 736
        ,  1.503    ,  3.094            // 737
        ,   1.68    ,  2.917            // 738
        ,   1.68    ,  3.094            // 739
        ,  1.503    ,  3.448            // 740
        ,  1.503    ,  3.271            // 741
        ,   1.68    ,  3.448            // 742
        ,   1.68    ,  3.271            // 743
        ,  2.033    ,  2.917            // 744
        ,  2.033    ,  3.094            // 745
        ,  1.856    ,  2.917            // 746
        ,  1.856    ,  3.094            // 747
        ,  2.033    ,  3.448            // 748
        ,  2.033    ,  3.271            // 749
        ,  1.856    ,  3.448            // 750
        ,  1.856    ,  3.271            // 751
        ,  1.503    ,  4.155            // 752
        ,  1.503    ,  3.978            // 753
        ,   1.68    ,  4.155            // 754
        ,   1.68    ,  3.978            // 755
        ,  1.503    ,  3.624            // 756
        ,  1.503    ,  3.801            // 757
        ,   1.68    ,  3.624            // 758
        ,   1.68    ,  3.801            // 759
        ,  2.033    ,  4.155            // 760
        ,  2.033    ,  3.978            // 761
        ,  1.856    ,  4.155            // 762
        ,  1.856    ,  3.978            // 763
        ,  2.033    ,  3.624            // 764
        ,  2.033    ,  3.801            // 765
        ,  1.856    ,  3.624            // 766
        ,  1.856    ,  3.801            // 767
        ,  0.088    ,  0.088            // 768
        ,  0.088    ,  0.265            // 769
        ,  0.265    ,  0.088            // 770
        ,  0.265    ,  0.265            // 771
        ,  0.088    ,  0.619            // 772
        ,  0.088    ,  0.442            // 773
        ,  0.265    ,  0.619            // 774
        ,  0.265    ,  0.442            // 775
        ,  0.619    ,  0.088            // 776
        ,  0.619    ,  0.265            // 777
        ,  0.442    ,  0.088            // 778
        ,  0.442    ,  0.265            // 779
        ,  0.619    ,  0.619            // 780
        ,  0.619    ,  0.442            // 781
        ,  0.442    ,  0.619            // 782
        ,  0.442    ,  0.442            // 783
        ,  0.088    ,  1.326            // 784
        ,  0.088    ,  1.149            // 785
        ,  0.265    ,  1.326            // 786
        ,  0.265    ,  1.149            // 787
        ,  0.088    ,  0.796            // 788
        ,  0.088    ,  0.972            // 789
        ,  0.265    ,  0.796            // 790
        ,  0.265    ,  0.972            // 791
        ,  0.619    ,  1.326            // 792
        ,  0.619    ,  1.149            // 793
        ,  0.442    ,  1.326            // 794
        ,  0.442    ,  1.149            // 795
        ,  0.619    ,  0.796            // 796
        ,  0.619    ,  0.972            // 797
        ,  0.442    ,  0.796            // 798
        ,  0.442    ,  0.972            // 799
        ,  1.326    ,  0.088            // 800
        ,  1.326    ,  0.265            // 801
        ,  1.149    ,  0.088            // 802
        ,  1.149    ,  0.265            // 803
        ,  1.326    ,  0.619            // 804
        ,  1.326    ,  0.442            // 805
        ,  1.149    ,  0.619            // 806
        ,  1.149    ,  0.442            // 807
        ,  0.796    ,  0.088            // 808
        ,  0.796    ,  0.265            // 809
        ,  0.972    ,  0.088            // 810
        ,  0.972    ,  0.265            // 811
        ,  0.796    ,  0.619            // 812
        ,  0.796    ,  0.442            // 813
        ,  0.972    ,  0.619            // 814
        ,  0.972    ,  0.442            // 815
        ,  1.326    ,  1.326            // 816
        ,  1.326    ,  1.149            // 817
        ,  1.149    ,  1.326            // 818
        ,  1.149    ,  1.149            // 819
        ,  1.326    ,  0.796            // 820
        ,  1.326    ,  0.972            // 821
        ,  1.149    ,  0.796            // 822
        ,  1.149    ,  0.972            // 823
        ,  0.796    ,  1.326            // 824
        ,  0.796    ,  1.149            // 825
        ,  0.972    ,  1.326            // 826
        ,  0.972    ,  1.149            // 827
        ,  0.796    ,  0.796            // 828
        ,  0.796    ,  0.972            // 829
        ,  0.972    ,  0.796            // 830
        ,  0.972    ,  0.972            // 831
        ,  0.088    ,   2.74            // 832
        ,  0.088    ,  2.564            // 833
        ,  0.265    ,   2.74            // 834
        ,  0.265    ,  2.564            // 835
        ,  0.088    ,   2.21            // 836
        ,  0.088    ,  2.387            // 837
        ,  0.265    ,   2.21            // 838
        ,  0.265    ,  2.387            // 839
        ,  0.619    ,   2.74            // 840
        ,  0.619    ,  2.564            // 841
        ,  0.442    ,   2.74            // 842
        ,  0.442    ,  2.564            // 843
        ,  0.619    ,   2.21            // 844
        ,  0.619    ,  2.387            // 845
        ,  0.442    ,   2.21            // 846
        ,  0.442    ,  2.387            // 847
        ,  0.088    ,  1.503            // 848
        ,  0.088    ,   1.68            // 849
        ,  0.265    ,  1.503            // 850
        ,  0.265    ,   1.68            // 851
        ,  0.088    ,  2.033            // 852
        ,  0.088    ,  1.856            // 853
        ,  0.265    ,  2.033            // 854
        ,  0.265    ,  1.856            // 855
        ,  0.619    ,  1.503            // 856
        ,  0.619    ,   1.68            // 857
        ,  0.442    ,  1.503            // 858
        ,  0.442    ,   1.68            // 859
        ,  0.619    ,  2.033            // 860
        ,  0.619    ,  1.856            // 861
        ,  0.442    ,  2.033            // 862
        ,  0.442    ,  1.856            // 863
        ,  1.326    ,   2.74            // 864
        ,  1.326    ,  2.564            // 865
        ,  1.149    ,   2.74            // 866
        ,  1.149    ,  2.564            // 867
        ,  1.326    ,   2.21            // 868
        ,  1.326    ,  2.387            // 869
        ,  1.149    ,   2.21            // 870
        ,  1.149    ,  2.387            // 871
        ,  0.796    ,   2.74            // 872
        ,  0.796    ,  2.564            // 873
        ,  0.972    ,   2.74            // 874
        ,  0.972    ,  2.564            // 875
        ,  0.796    ,   2.21            // 876
        ,  0.796    ,  2.387            // 877
        ,  0.972    ,   2.21            // 878
        ,  0.972    ,  2.387            // 879
        ,  1.326    ,  1.503            // 880
        ,  1.326    ,   1.68            // 881
        ,  1.149    ,  1.503            // 882
        ,  1.149    ,   1.68            // 883
        ,  1.326    ,  2.033            // 884
        ,  1.326    ,  1.856            // 885
        ,  1.149    ,  2.033            // 886
        ,  1.149    ,  1.856            // 887
        ,  0.796    ,  1.503            // 888
        ,  0.796    ,   1.68            // 889
        ,  0.972    ,  1.503            // 890
        ,  0.972    ,   1.68            // 891
        ,  0.796    ,  2.033            // 892
        ,  0.796    ,  1.856            // 893
        ,  0.972    ,  2.033            // 894
        ,  0.972    ,  1.856            // 895
        ,   2.74    ,  0.088            // 896
        ,   2.74    ,  0.265            // 897
        ,  2.564    ,  0.088            // 898
        ,  2.564    ,  0.265            // 899
        ,   2.74    ,  0.619            // 900
        ,   2.74    ,  0.442            // 901
        ,  2.564    ,  0.619            // 902
        ,  2.564    ,  0.442            // 903
        ,   2.21    ,  0.088            // 904
        ,   2.21    ,  0.265            // 905
        ,  2.387    ,  0.088            // 906
        ,  2.387    ,  0.265            // 907
        ,   2.21    ,  0.619            // 908
        ,   2.21    ,  0.442            // 909
        ,  2.387    ,  0.619            // 910
        ,  2.387    ,  0.442            // 911
        ,   2.74    ,  1.326            // 912
        ,   2.74    ,  1.149            // 913
        ,  2.564    ,  1.326            // 914
        ,  2.564    ,  1.149            // 915
        ,   2.74    ,  0.796            // 916
        ,   2.74    ,  0.972            // 917
        ,  2.564    ,  0.796            // 918
        ,  2.564    ,  0.972            // 919
        ,   2.21    ,  1.326            // 920
        ,   2.21    ,  1.149            // 921
        ,  2.387    ,  1.326            // 922
        ,  2.387    ,  1.149            // 923
        ,   2.21    ,  0.796            // 924
        ,   2.21    ,  0.972            // 925
        ,  2.387    ,  0.796            // 926
        ,  2.387    ,  0.972            // 927
        ,  1.503    ,  0.088            // 928
        ,  1.503    ,  0.265            // 929
        ,   1.68    ,  0.088            // 930
        ,   1.68    ,  0.265            // 931
        ,  1.503    ,  0.619            // 932
        ,  1.503    ,  0.442            // 933
        ,   1.68    ,  0.619            // 934
        ,   1.68    ,  0.442            // 935
        ,  2.033    ,  0.088            // 936
        ,  2.033    ,  0.265            // 937
        ,  1.856    ,  0.088            // 938
        ,  1.856    ,  0.265            // 939
        ,  2.033    ,  0.619            // 940
        ,  2.033    ,  0.442            // 941
        ,  1.856    ,  0.619            // 942
        ,  1.856    ,  0.442            // 943
        ,  1.503    ,  1.326            // 944
        ,  1.503    ,  1.149            // 945
        ,   1.68    ,  1.326            // 946
        ,   1.68    ,  1.149            // 947
        ,  1.503    ,  0.796            // 948
        ,  1.503    ,  0.972            // 949
        ,   1.68    ,  0.796            // 950
        ,   1.68    ,  0.972            // 951
        ,  2.033    ,  1.326            // 952
        ,  2.033    ,  1.149            // 953
        ,  1.856    ,  1.326            // 954
        ,  1.856    ,  1.149            // 955
        ,  2.033    ,  0.796            // 956
        ,  2.033    ,  0.972            // 957
        ,  1.856    ,  0.796            // 958
        ,  1.856    ,  0.972            // 959
        ,   2.74    ,   2.74            // 960
        ,   2.74    ,  2.564            // 961
        ,  2.564    ,   2.74            // 962
        ,  2.564    ,  2.564            // 963
        ,   2.74    ,   2.21            // 964
        ,   2.74    ,  2.387            // 965
        ,  2.564    ,   2.21            // 966
        ,  2.564    ,  2.387            // 967
        ,   2.21    ,   2.74            // 968
        ,   2.21    ,  2.564            // 969
        ,  2.387    ,   2.74            // 970
        ,  2.387    ,  2.564            // 971
        ,   2.21    ,   2.21            // 972
        ,   2.21    ,  2.387            // 973
        ,  2.387    ,   2.21            // 974
        ,  2.387    ,  2.387            // 975
        ,   2.74    ,  1.503            // 976
        ,   2.74    ,   1.68            // 977
        ,  2.564    ,  1.503            // 978
        ,  2.564    ,   1.68            // 979
        ,   2.74    ,  2.033            // 980
        ,   2.74    ,  1.856            // 981
        ,  2.564    ,  2.033            // 982
        ,  2.564    ,  1.856            // 983
        ,   2.21    ,  1.503            // 984
        ,   2.21    ,   1.68            // 985
        ,  2.387    ,  1.503            // 986
        ,  2.387    ,   1.68            // 987
        ,   2.21    ,  2.033            // 988
        ,   2.21    ,  1.856            // 989
        ,  2.387    ,  2.033            // 990
        ,  2.387    ,  1.856            // 991
        ,  1.503    ,   2.74            // 992
        ,  1.503    ,  2.564            // 993
        ,   1.68    ,   2.74            // 994
        ,   1.68    ,  2.564            // 995
        ,  1.503    ,   2.21            // 996
        ,  1.503    ,  2.387            // 997
        ,   1.68    ,   2.21            // 998
        ,   1.68    ,  2.387            // 999
        ,  2.033    ,   2.74            // 1000
        ,  2.033    ,  2.564            // 1001
        ,  1.856    ,   2.74            // 1002
        ,  1.856    ,  2.564            // 1003
        ,  2.033    ,   2.21            // 1004
        ,  2.033    ,  2.387            // 1005
        ,  1.856    ,   2.21            // 1006
        ,  1.856    ,  2.387            // 1007
        ,  1.503    ,  1.503            // 1008
        ,  1.503    ,   1.68            // 1009
        ,   1.68    ,  1.503            // 1010
        ,   1.68    ,   1.68            // 1011
        ,  1.503    ,  2.033            // 1012
        ,  1.503    ,  1.856            // 1013
        ,   1.68    ,  2.033            // 1014
        ,   1.68    ,  1.856            // 1015
        ,  2.033    ,  1.503            // 1016
        ,  2.033    ,   1.68            // 1017
        ,  1.856    ,  1.503            // 1018
        ,  1.856    ,   1.68            // 1019
        ,  2.033    ,  2.033            // 1020
        ,  2.033    ,  1.856            // 1021
        ,  1.856    ,  2.033            // 1022
        ,  1.856    ,  1.856            // 1023
        ,  5.569    , -5.569            // 1024
        ,  5.569    , -5.392            // 1025
        ,  5.392    , -5.569            // 1026
        ,  5.392    , -5.392            // 1027
        ,  5.569    , -5.039            // 1028
        ,  5.569    , -5.216            // 1029
        ,  5.392    , -5.039            // 1030
        ,  5.392    , -5.216            // 1031
        ,  5.039    , -5.569            // 1032
        ,  5.039    , -5.392            // 1033
        ,  5.216    , -5.569            // 1034
        ,  5.216    , -5.392            // 1035
        ,  5.039    , -5.039            // 1036
        ,  5.039    , -5.216            // 1037
        ,  5.216    , -5.039            // 1038
        ,  5.216    , -5.216            // 1039
        ,  5.569    , -4.332            // 1040
        ,  5.569    , -4.508            // 1041
        ,  5.392    , -4.332            // 1042
        ,  5.392    , -4.508            // 1043
        ,  5.569    , -4.862            // 1044
        ,  5.569    , -4.685            // 1045
        ,  5.392    , -4.862            // 1046
        ,  5.392    , -4.685            // 1047
        ,  5.039    , -4.332            // 1048
        ,  5.039    , -4.508            // 1049
        ,  5.216    , -4.332            // 1050
        ,  5.216    , -4.508            // 1051
        ,  5.039    , -4.862            // 1052
        ,  5.039    , -4.685            // 1053
        ,  5.216    , -4.862            // 1054
        ,  5.216    , -4.685            // 1055
        ,  4.332    , -5.569            // 1056
        ,  4.332    , -5.392            // 1057
        ,  4.508    , -5.569            // 1058
        ,  4.508    , -5.392            // 1059
        ,  4.332    , -5.039            // 1060
        ,  4.332    , -5.216            // 1061
        ,  4.508    , -5.039            // 1062
        ,  4.508    , -5.216            // 1063
        ,  4.862    , -5.569            // 1064
        ,  4.862    , -5.392            // 1065
        ,  4.685    , -5.569            // 1066
        ,  4.685    , -5.392            // 1067
        ,  4.862    , -5.039            // 1068
        ,  4.862    , -5.216            // 1069
        ,  4.685    , -5.039            // 1070
        ,  4.685    , -5.216            // 1071
        ,  4.332    , -4.332            // 1072
        ,  4.332    , -4.508            // 1073
        ,  4.508    , -4.332            // 1074
        ,  4.508    , -4.508            // 1075
        ,  4.332    , -4.862            // 1076
        ,  4.332    , -4.685            // 1077
        ,  4.508    , -4.862            // 1078
        ,  4.508    , -4.685            // 1079
        ,  4.862    , -4.332            // 1080
        ,  4.862    , -4.508            // 1081
        ,  4.685    , -4.332            // 1082
        ,  4.685    , -4.508            // 1083
        ,  4.862    , -4.862            // 1084
        ,  4.862    , -4.685            // 1085
        ,  4.685    , -4.862            // 1086
        ,  4.685    , -4.685            // 1087
        ,  5.569    , -2.917            // 1088
        ,  5.569    , -3.094            // 1089
        ,  5.392    , -2.917            // 1090
        ,  5.392    , -3.094            // 1091
        ,  5.569    , -3.448            // 1092
        ,  5.569    , -3.271            // 1093
        ,  5.392    , -3.448            // 1094
        ,  5.392    , -3.271            // 1095
        ,  5.039    , -2.917            // 1096
        ,  5.039    , -3.094            // 1097
        ,  5.216    , -2.917            // 1098
        ,  5.216    , -3.094            // 1099
        ,  5.039    , -3.448            // 1100
        ,  5.039    , -3.271            // 1101
        ,  5.216    , -3.448            // 1102
        ,  5.216    , -3.271            // 1103
        ,  5.569    , -4.155            // 1104
        ,  5.569    , -3.978            // 1105
        ,  5.392    , -4.155            // 1106
        ,  5.392    , -3.978            // 1107
        ,  5.569    , -3.624            // 1108
        ,  5.569    , -3.801            // 1109
        ,  5.392    , -3.624            // 1110
        ,  5.392    , -3.801            // 1111
        ,  5.039    , -4.155            // 1112
        ,  5.039    , -3.978            // 1113
        ,  5.216    , -4.155            // 1114
        ,  5.216    , -3.978            // 1115
        ,  5.039    , -3.624            // 1116
        ,  5.039    , -3.801            // 1117
        ,  5.216    , -3.624            // 1118
        ,  5.216    , -3.801            // 1119
        ,  4.332    , -2.917            // 1120
        ,  4.332    , -3.094            // 1121
        ,  4.508    , -2.917            // 1122
        ,  4.508    , -3.094            // 1123
        ,  4.332    , -3.448            // 1124
        ,  4.332    , -3.271            // 1125
        ,  4.508    , -3.448            // 1126
        ,  4.508    , -3.271            // 1127
        ,  4.862    , -2.917            // 1128
        ,  4.862    , -3.094            // 1129
        ,  4.685    , -2.917            // 1130
        ,  4.685    , -3.094            // 1131
        ,  4.862    , -3.448            // 1132
        ,  4.862    , -3.271            // 1133
        ,  4.685    , -3.448            // 1134
        ,  4.685    , -3.271            // 1135
        ,  4.332    , -4.155            // 1136
        ,  4.332    , -3.978            // 1137
        ,  4.508    , -4.155            // 1138
        ,  4.508    , -3.978            // 1139
        ,  4.332    , -3.624            // 1140
        ,  4.332    , -3.801            // 1141
        ,  4.508    , -3.624            // 1142
        ,  4.508    , -3.801            // 1143
        ,  4.862    , -4.155            // 1144
        ,  4.862    , -3.978            // 1145
        ,  4.685    , -4.155            // 1146
        ,  4.685    , -3.978            // 1147
        ,  4.862    , -3.624            // 1148
        ,  4.862    , -3.801            // 1149
        ,  4.685    , -3.624            // 1150
        ,  4.685    , -3.801            // 1151
        ,  2.917    , -5.569            // 1152
        ,  2.917    , -5.392            // 1153
        ,  3.094    , -5.569            // 1154
        ,  3.094    , -5.392            // 1155
        ,  2.917    , -5.039            // 1156
        ,  2.917    , -5.216            // 1157
        ,  3.094    , -5.039            // 1158
        ,  3.094    , -5.216            // 1159
        ,  3.448    , -5.569            // 1160
        ,  3.448    , -5.392            // 1161
        ,  3.271    , -5.569            // 1162
        ,  3.271    , -5.392            // 1163
        ,  3.448    , -5.039            // 1164
        ,  3.448    , -5.216            // 1165
        ,  3.271    , -5.039            // 1166
        ,  3.271    , -5.216            // 1167
        ,  2.917    , -4.332            // 1168
        ,  2.917    , -4.508            // 1169
        ,  3.094    , -4.332            // 1170
        ,  3.094    , -4.508            // 1171
        ,  2.917    , -4.862            // 1172
        ,  2.917    , -4.685            // 1173
        ,  3.094    , -4.862            // 1174
        ,  3.094    , -4.685            // 1175
        ,  3.448    , -4.332            // 1176
        ,  3.448    , -4.508            // 1177
        ,  3.271    , -4.332            // 1178
        ,  3.271    , -4.508            // 1179
        ,  3.448    , -4.862            // 1180
        ,  3.448    , -4.685            // 1181
        ,  3.271    , -4.862            // 1182
        ,  3.271    , -4.685            // 1183
        ,  4.155    , -5.569            // 1184
        ,  4.155    , -5.392            // 1185
        ,  3.978    , -5.569            // 1186
        ,  3.978    , -5.392            // 1187
        ,  4.155    , -5.039            // 1188
        ,  4.155    , -5.216            // 1189
        ,  3.978    , -5.039            // 1190
        ,  3.978    , -5.216            // 1191
        ,  3.624    , -5.569            // 1192
        ,  3.624    , -5.392            // 1193
        ,  3.801    , -5.569            // 1194
        ,  3.801    , -5.392            // 1195
        ,  3.624    , -5.039            // 1196
        ,  3.624    , -5.216            // 1197
        ,  3.801    , -5.039            // 1198
        ,  3.801    , -5.216            // 1199
        ,  4.155    , -4.332            // 1200
        ,  4.155    , -4.508            // 1201
        ,  3.978    , -4.332            // 1202
        ,  3.978    , -4.508            // 1203
        ,  4.155    , -4.862            // 1204
        ,  4.155    , -4.685            // 1205
        ,  3.978    , -4.862            // 1206
        ,  3.978    , -4.685            // 1207
        ,  3.624    , -4.332            // 1208
        ,  3.624    , -4.508            // 1209
        ,  3.801    , -4.332            // 1210
        ,  3.801    , -4.508            // 1211
        ,  3.624    , -4.862            // 1212
        ,  3.624    , -4.685            // 1213
        ,  3.801    , -4.862            // 1214
        ,  3.801    , -4.685            // 1215
        ,  2.917    , -2.917            // 1216
        ,  2.917    , -3.094            // 1217
        ,  3.094    , -2.917            // 1218
        ,  3.094    , -3.094            // 1219
        ,  2.917    , -3.448            // 1220
        ,  2.917    , -3.271            // 1221
        ,  3.094    , -3.448            // 1222
        ,  3.094    , -3.271            // 1223
        ,  3.448    , -2.917            // 1224
        ,  3.448    , -3.094            // 1225
        ,  3.271    , -2.917            // 1226
        ,  3.271    , -3.094            // 1227
        ,  3.448    , -3.448            // 1228
        ,  3.448    , -3.271            // 1229
        ,  3.271    , -3.448            // 1230
        ,  3.271    , -3.271            // 1231
        ,  2.917    , -4.155            // 1232
        ,  2.917    , -3.978            // 1233
        ,  3.094    , -4.155            // 1234
        ,  3.094    , -3.978            // 1235
        ,  2.917    , -3.624            // 1236
        ,  2.917    , -3.801            // 1237
        ,  3.094    , -3.624            // 1238
        ,  3.094    , -3.801            // 1239
        ,  3.448    , -4.155            // 1240
        ,  3.448    , -3.978            // 1241
        ,  3.271    , -4.155            // 1242
        ,  3.271    , -3.978            // 1243
        ,  3.448    , -3.624            // 1244
        ,  3.448    , -3.801            // 1245
        ,  3.271    , -3.624            // 1246
        ,  3.271    , -3.801            // 1247
        ,  4.155    , -2.917            // 1248
        ,  4.155    , -3.094            // 1249
        ,  3.978    , -2.917            // 1250
        ,  3.978    , -3.094            // 1251
        ,  4.155    , -3.448            // 1252
        ,  4.155    , -3.271            // 1253
        ,  3.978    , -3.448            // 1254
        ,  3.978    , -3.271            // 1255
        ,  3.624    , -2.917            // 1256
        ,  3.624    , -3.094            // 1257
        ,  3.801    , -2.917            // 1258
        ,  3.801    , -3.094            // 1259
        ,  3.624    , -3.448            // 1260
        ,  3.624    , -3.271            // 1261
        ,  3.801    , -3.448            // 1262
        ,  3.801    , -3.271            // 1263
        ,  4.155    , -4.155            // 1264
        ,  4.155    , -3.978            // 1265
        ,  3.978    , -4.155            // 1266
        ,  3.978    , -3.978            // 1267
        ,  4.155    , -3.624            // 1268
        ,  4.155    , -3.801            // 1269
        ,  3.978    , -3.624            // 1270
        ,  3.978    , -3.801            // 1271
        ,  3.624    , -4.155            // 1272
        ,  3.624    , -3.978            // 1273
        ,  3.801    , -4.155            // 1274
        ,  3.801    , -3.978            // 1275
        ,  3.624    , -3.624            // 1276
        ,  3.624    , -3.801            // 1277
        ,  3.801    , -3.624            // 1278
        ,  3.801    , -3.801            // 1279
        ,  5.569    , -0.088            // 1280
        ,  5.569    , -0.265            // 1281
        ,  5.392    , -0.088            // 1282
        ,  5.392    , -0.265            // 1283
        ,  5.569    , -0.619            // 1284
        ,  5.569    , -0.442            // 1285
        ,  5.392    , -0.619            // 1286
        ,  5.392    , -0.442            // 1287
        ,  5.039    , -0.088            // 1288
        ,  5.039    , -0.265            // 1289
        ,  5.216    , -0.088            // 1290
        ,  5.216    , -0.265            // 1291
        ,  5.039    , -0.619            // 1292
        ,  5.039    , -0.442            // 1293
        ,  5.216    , -0.619            // 1294
        ,  5.216    , -0.442            // 1295
        ,  5.569    , -1.326            // 1296
        ,  5.569    , -1.149            // 1297
        ,  5.392    , -1.326            // 1298
        ,  5.392    , -1.149            // 1299
        ,  5.569    , -0.796            // 1300
        ,  5.569    , -0.972            // 1301
        ,  5.392    , -0.796            // 1302
        ,  5.392    , -0.972            // 1303
        ,  5.039    , -1.326            // 1304
        ,  5.039    , -1.149            // 1305
        ,  5.216    , -1.326            // 1306
        ,  5.216    , -1.149            // 1307
        ,  5.039    , -0.796            // 1308
        ,  5.039    , -0.972            // 1309
        ,  5.216    , -0.796            // 1310
        ,  5.216    , -0.972            // 1311
        ,  4.332    , -0.088            // 1312
        ,  4.332    , -0.265            // 1313
        ,  4.508    , -0.088            // 1314
        ,  4.508    , -0.265            // 1315
        ,  4.332    , -0.619            // 1316
        ,  4.332    , -0.442            // 1317
        ,  4.508    , -0.619            // 1318
        ,  4.508    , -0.442            // 1319
        ,  4.862    , -0.088            // 1320
        ,  4.862    , -0.265            // 1321
        ,  4.685    , -0.088            // 1322
        ,  4.685    , -0.265            // 1323
        ,  4.862    , -0.619            // 1324
        ,  4.862    , -0.442            // 1325
        ,  4.685    , -0.619            // 1326
        ,  4.685    , -0.442            // 1327
        ,  4.332    , -1.326            // 1328
        ,  4.332    , -1.149            // 1329
        ,  4.508    , -1.326            // 1330
        ,  4.508    , -1.149            // 1331
        ,  4.332    , -0.796            // 1332
        ,  4.332    , -0.972            // 1333
        ,  4.508    , -0.796            // 1334
        ,  4.508    , -0.972            // 1335
        ,  4.862    , -1.326            // 1336
        ,  4.862    , -1.149            // 1337
        ,  4.685    , -1.326            // 1338
        ,  4.685    , -1.149            // 1339
        ,  4.862    , -0.796            // 1340
        ,  4.862    , -0.972            // 1341
        ,  4.685    , -0.796            // 1342
        ,  4.685    , -0.972            // 1343
        ,  5.569    ,  -2.74            // 1344
        ,  5.569    , -2.564            // 1345
        ,  5.392    ,  -2.74            // 1346
        ,  5.392    , -2.564            // 1347
        ,  5.569    ,  -2.21            // 1348
        ,  5.569    , -2.387            // 1349
        ,  5.392    ,  -2.21            // 1350
        ,  5.392    , -2.387            // 1351
        ,  5.039    ,  -2.74            // 1352
        ,  5.039    , -2.564            // 1353
        ,  5.216    ,  -2.74            // 1354
        ,  5.216    , -2.564            // 1355
        ,  5.039    ,  -2.21            // 1356
        ,  5.039    , -2.387            // 1357
        ,  5.216    ,  -2.21            // 1358
        ,  5.216    , -2.387            // 1359
        ,  5.569    , -1.503            // 1360
        ,  5.569    ,  -1.68            // 1361
        ,  5.392    , -1.503            // 1362
        ,  5.392    ,  -1.68            // 1363
        ,  5.569    , -2.033            // 1364
        ,  5.569    , -1.856            // 1365
        ,  5.392    , -2.033            // 1366
        ,  5.392    , -1.856            // 1367
        ,  5.039    , -1.503            // 1368
        ,  5.039    ,  -1.68            // 1369
        ,  5.216    , -1.503            // 1370
        ,  5.216    ,  -1.68            // 1371
        ,  5.039    , -2.033            // 1372
        ,  5.039    , -1.856            // 1373
        ,  5.216    , -2.033            // 1374
        ,  5.216    , -1.856            // 1375
        ,  4.332    ,  -2.74            // 1376
        ,  4.332    , -2.564            // 1377
        ,  4.508    ,  -2.74            // 1378
        ,  4.508    , -2.564            // 1379
        ,  4.332    ,  -2.21            // 1380
        ,  4.332    , -2.387            // 1381
        ,  4.508    ,  -2.21            // 1382
        ,  4.508    , -2.387            // 1383
        ,  4.862    ,  -2.74            // 1384
        ,  4.862    , -2.564            // 1385
        ,  4.685    ,  -2.74            // 1386
        ,  4.685    , -2.564            // 1387
        ,  4.862    ,  -2.21            // 1388
        ,  4.862    , -2.387            // 1389
        ,  4.685    ,  -2.21            // 1390
        ,  4.685    , -2.387            // 1391
        ,  4.332    , -1.503            // 1392
        ,  4.332    ,  -1.68            // 1393
        ,  4.508    , -1.503            // 1394
        ,  4.508    ,  -1.68            // 1395
        ,  4.332    , -2.033            // 1396
        ,  4.332    , -1.856            // 1397
        ,  4.508    , -2.033            // 1398
        ,  4.508    , -1.856            // 1399
        ,  4.862    , -1.503            // 1400
        ,  4.862    ,  -1.68            // 1401
        ,  4.685    , -1.503            // 1402
        ,  4.685    ,  -1.68            // 1403
        ,  4.862    , -2.033            // 1404
        ,  4.862    , -1.856            // 1405
        ,  4.685    , -2.033            // 1406
        ,  4.685    , -1.856            // 1407
        ,  2.917    , -0.088            // 1408
        ,  2.917    , -0.265            // 1409
        ,  3.094    , -0.088            // 1410
        ,  3.094    , -0.265            // 1411
        ,  2.917    , -0.619            // 1412
        ,  2.917    , -0.442            // 1413
        ,  3.094    , -0.619            // 1414
        ,  3.094    , -0.442            // 1415
        ,  3.448    , -0.088            // 1416
        ,  3.448    , -0.265            // 1417
        ,  3.271    , -0.088            // 1418
        ,  3.271    , -0.265            // 1419
        ,  3.448    , -0.619            // 1420
        ,  3.448    , -0.442            // 1421
        ,  3.271    , -0.619            // 1422
        ,  3.271    , -0.442            // 1423
        ,  2.917    , -1.326            // 1424
        ,  2.917    , -1.149            // 1425
        ,  3.094    , -1.326            // 1426
        ,  3.094    , -1.149            // 1427
        ,  2.917    , -0.796            // 1428
        ,  2.917    , -0.972            // 1429
        ,  3.094    , -0.796            // 1430
        ,  3.094    , -0.972            // 1431
        ,  3.448    , -1.326            // 1432
        ,  3.448    , -1.149            // 1433
        ,  3.271    , -1.326            // 1434
        ,  3.271    , -1.149            // 1435
        ,  3.448    , -0.796            // 1436
        ,  3.448    , -0.972            // 1437
        ,  3.271    , -0.796            // 1438
        ,  3.271    , -0.972            // 1439
        ,  4.155    , -0.088            // 1440
        ,  4.155    , -0.265            // 1441
        ,  3.978    , -0.088            // 1442
        ,  3.978    , -0.265            // 1443
        ,  4.155    , -0.619            // 1444
        ,  4.155    , -0.442            // 1445
        ,  3.978    , -0.619            // 1446
        ,  3.978    , -0.442            // 1447
        ,  3.624    , -0.088            // 1448
        ,  3.624    , -0.265            // 1449
        ,  3.801    , -0.088            // 1450
        ,  3.801    , -0.265            // 1451
        ,  3.624    , -0.619            // 1452
        ,  3.624    , -0.442            // 1453
        ,  3.801    , -0.619            // 1454
        ,  3.801    , -0.442            // 1455
        ,  4.155    , -1.326            // 1456
        ,  4.155    , -1.149            // 1457
        ,  3.978    , -1.326            // 1458
        ,  3.978    , -1.149            // 1459
        ,  4.155    , -0.796            // 1460
        ,  4.155    , -0.972            // 1461
        ,  3.978    , -0.796            // 1462
        ,  3.978    , -0.972            // 1463
        ,  3.624    , -1.326            // 1464
        ,  3.624    , -1.149            // 1465
        ,  3.801    , -1.326            // 1466
        ,  3.801    , -1.149            // 1467
        ,  3.624    , -0.796            // 1468
        ,  3.624    , -0.972            // 1469
        ,  3.801    , -0.796            // 1470
        ,  3.801    , -0.972            // 1471
        ,  2.917    ,  -2.74            // 1472
        ,  2.917    , -2.564            // 1473
        ,  3.094    ,  -2.74            // 1474
        ,  3.094    , -2.564            // 1475
        ,  2.917    ,  -2.21            // 1476
        ,  2.917    , -2.387            // 1477
        ,  3.094    ,  -2.21            // 1478
        ,  3.094    , -2.387            // 1479
        ,  3.448    ,  -2.74            // 1480
        ,  3.448    , -2.564            // 1481
        ,  3.271    ,  -2.74            // 1482
        ,  3.271    , -2.564            // 1483
        ,  3.448    ,  -2.21            // 1484
        ,  3.448    , -2.387            // 1485
        ,  3.271    ,  -2.21            // 1486
        ,  3.271    , -2.387            // 1487
        ,  2.917    , -1.503            // 1488
        ,  2.917    ,  -1.68            // 1489
        ,  3.094    , -1.503            // 1490
        ,  3.094    ,  -1.68            // 1491
        ,  2.917    , -2.033            // 1492
        ,  2.917    , -1.856            // 1493
        ,  3.094    , -2.033            // 1494
        ,  3.094    , -1.856            // 1495
        ,  3.448    , -1.503            // 1496
        ,  3.448    ,  -1.68            // 1497
        ,  3.271    , -1.503            // 1498
        ,  3.271    ,  -1.68            // 1499
        ,  3.448    , -2.033            // 1500
        ,  3.448    , -1.856            // 1501
        ,  3.271    , -2.033            // 1502
        ,  3.271    , -1.856            // 1503
        ,  4.155    ,  -2.74            // 1504
        ,  4.155    , -2.564            // 1505
        ,  3.978    ,  -2.74            // 1506
        ,  3.978    , -2.564            // 1507
        ,  4.155    ,  -2.21            // 1508
        ,  4.155    , -2.387            // 1509
        ,  3.978    ,  -2.21            // 1510
        ,  3.978    , -2.387            // 1511
        ,  3.624    ,  -2.74            // 1512
        ,  3.624    , -2.564            // 1513
        ,  3.801    ,  -2.74            // 1514
        ,  3.801    , -2.564            // 1515
        ,  3.624    ,  -2.21            // 1516
        ,  3.624    , -2.387            // 1517
        ,  3.801    ,  -2.21            // 1518
        ,  3.801    , -2.387            // 1519
        ,  4.155    , -1.503            // 1520
        ,  4.155    ,  -1.68            // 1521
        ,  3.978    , -1.503            // 1522
        ,  3.978    ,  -1.68            // 1523
        ,  4.155    , -2.033            // 1524
        ,  4.155    , -1.856            // 1525
        ,  3.978    , -2.033            // 1526
        ,  3.978    , -1.856            // 1527
        ,  3.624    , -1.503            // 1528
        ,  3.624    ,  -1.68            // 1529
        ,  3.801    , -1.503            // 1530
        ,  3.801    ,  -1.68            // 1531
        ,  3.624    , -2.033            // 1532
        ,  3.624    , -1.856            // 1533
        ,  3.801    , -2.033            // 1534
        ,  3.801    , -1.856            // 1535
        ,  0.088    , -5.569            // 1536
        ,  0.088    , -5.392            // 1537
        ,  0.265    , -5.569            // 1538
        ,  0.265    , -5.392            // 1539
        ,  0.088    , -5.039            // 1540
        ,  0.088    , -5.216            // 1541
        ,  0.265    , -5.039            // 1542
        ,  0.265    , -5.216            // 1543
        ,  0.619    , -5.569            // 1544
        ,  0.619    , -5.392            // 1545
        ,  0.442    , -5.569            // 1546
        ,  0.442    , -5.392            // 1547
        ,  0.619    , -5.039            // 1548
        ,  0.619    , -5.216            // 1549
        ,  0.442    , -5.039            // 1550
        ,  0.442    , -5.216            // 1551
        ,  0.088    , -4.332            // 1552
        ,  0.088    , -4.508            // 1553
        ,  0.265    , -4.332            // 1554
        ,  0.265    , -4.508            // 1555
        ,  0.088    , -4.862            // 1556
        ,  0.088    , -4.685            // 1557
        ,  0.265    , -4.862            // 1558
        ,  0.265    , -4.685            // 1559
        ,  0.619    , -4.332            // 1560
        ,  0.619    , -4.508            // 1561
        ,  0.442    , -4.332            // 1562
        ,  0.442    , -4.508            // 1563
        ,  0.619    , -4.862            // 1564
        ,  0.619    , -4.685            // 1565
        ,  0.442    , -4.862            // 1566
        ,  0.442    , -4.685            // 1567
        ,  1.326    , -5.569            // 1568
        ,  1.326    , -5.392            // 1569
        ,  1.149    , -5.569            // 1570
        ,  1.149    , -5.392            // 1571
        ,  1.326    , -5.039            // 1572
        ,  1.326    , -5.216            // 1573
        ,  1.149    , -5.039            // 1574
        ,  1.149    , -5.216            // 1575
        ,  0.796    , -5.569            // 1576
        ,  0.796    , -5.392            // 1577
        ,  0.972    , -5.569            // 1578
        ,  0.972    , -5.392            // 1579
        ,  0.796    , -5.039            // 1580
        ,  0.796    , -5.216            // 1581
        ,  0.972    , -5.039            // 1582
        ,  0.972    , -5.216            // 1583
        ,  1.326    , -4.332            // 1584
        ,  1.326    , -4.508            // 1585
        ,  1.149    , -4.332            // 1586
        ,  1.149    , -4.508            // 1587
        ,  1.326    , -4.862            // 1588
        ,  1.326    , -4.685            // 1589
        ,  1.149    , -4.862            // 1590
        ,  1.149    , -4.685            // 1591
        ,  0.796    , -4.332            // 1592
        ,  0.796    , -4.508            // 1593
        ,  0.972    , -4.332            // 1594
        ,  0.972    , -4.508            // 1595
        ,  0.796    , -4.862            // 1596
        ,  0.796    , -4.685            // 1597
        ,  0.972    , -4.862            // 1598
        ,  0.972    , -4.685            // 1599
        ,  0.088    , -2.917            // 1600
        ,  0.088    , -3.094            // 1601
        ,  0.265    , -2.917            // 1602
        ,  0.265    , -3.094            // 1603
        ,  0.088    , -3.448            // 1604
        ,  0.088    , -3.271            // 1605
        ,  0.265    , -3.448            // 1606
        ,  0.265    , -3.271            // 1607
        ,  0.619    , -2.917            // 1608
        ,  0.619    , -3.094            // 1609
        ,  0.442    , -2.917            // 1610
        ,  0.442    , -3.094            // 1611
        ,  0.619    , -3.448            // 1612
        ,  0.619    , -3.271            // 1613
        ,  0.442    , -3.448            // 1614
        ,  0.442    , -3.271            // 1615
        ,  0.088    , -4.155            // 1616
        ,  0.088    , -3.978            // 1617
        ,  0.265    , -4.155            // 1618
        ,  0.265    , -3.978            // 1619
        ,  0.088    , -3.624            // 1620
        ,  0.088    , -3.801            // 1621
        ,  0.265    , -3.624            // 1622
        ,  0.265    , -3.801            // 1623
        ,  0.619    , -4.155            // 1624
        ,  0.619    , -3.978            // 1625
        ,  0.442    , -4.155            // 1626
        ,  0.442    , -3.978            // 1627
        ,  0.619    , -3.624            // 1628
        ,  0.619    , -3.801            // 1629
        ,  0.442    , -3.624            // 1630
        ,  0.442    , -3.801            // 1631
        ,  1.326    , -2.917            // 1632
        ,  1.326    , -3.094            // 1633
        ,  1.149    , -2.917            // 1634
        ,  1.149    , -3.094            // 1635
        ,  1.326    , -3.448            // 1636
        ,  1.326    , -3.271            // 1637
        ,  1.149    , -3.448            // 1638
        ,  1.149    , -3.271            // 1639
        ,  0.796    , -2.917            // 1640
        ,  0.796    , -3.094            // 1641
        ,  0.972    , -2.917            // 1642
        ,  0.972    , -3.094            // 1643
        ,  0.796    , -3.448            // 1644
        ,  0.796    , -3.271            // 1645
        ,  0.972    , -3.448            // 1646
        ,  0.972    , -3.271            // 1647
        ,  1.326    , -4.155            // 1648
        ,  1.326    , -3.978            // 1649
        ,  1.149    , -4.155            // 1650
        ,  1.149    , -3.978            // 1651
        ,  1.326    , -3.624            // 1652
        ,  1.326    , -3.801            // 1653
        ,  1.149    , -3.624            // 1654
        ,  1.149    , -3.801            // 1655
        ,  0.796    , -4.155            // 1656
        ,  0.796    , -3.978            // 1657
        ,  0.972    , -4.155            // 1658
        ,  0.972    , -3.978            // 1659
        ,  0.796    , -3.624            // 1660
        ,  0.796    , -3.801            // 1661
        ,  0.972    , -3.624            // 1662
        ,  0.972    , -3.801            // 1663
        ,   2.74    , -5.569            // 1664
        ,   2.74    , -5.392            // 1665
        ,  2.564    , -5.569            // 1666
        ,  2.564    , -5.392            // 1667
        ,   2.74    , -5.039            // 1668
        ,   2.74    , -5.216            // 1669
        ,  2.564    , -5.039            // 1670
        ,  2.564    , -5.216            // 1671
        ,   2.21    , -5.569            // 1672
        ,   2.21    , -5.392            // 1673
        ,  2.387    , -5.569            // 1674
        ,  2.387    , -5.392            // 1675
        ,   2.21    , -5.039            // 1676
        ,   2.21    , -5.216            // 1677
        ,  2.387    , -5.039            // 1678
        ,  2.387    , -5.216            // 1679
        ,   2.74    , -4.332            // 1680
        ,   2.74    , -4.508            // 1681
        ,  2.564    , -4.332            // 1682
        ,  2.564    , -4.508            // 1683
        ,   2.74    , -4.862            // 1684
        ,   2.74    , -4.685            // 1685
        ,  2.564    , -4.862            // 1686
        ,  2.564    , -4.685            // 1687
        ,   2.21    , -4.332            // 1688
        ,   2.21    , -4.508            // 1689
        ,  2.387    , -4.332            // 1690
        ,  2.387    , -4.508            // 1691
        ,   2.21    , -4.862            // 1692
        ,   2.21    , -4.685            // 1693
        ,  2.387    , -4.862            // 1694
        ,  2.387    , -4.685            // 1695
        ,  1.503    , -5.569            // 1696
        ,  1.503    , -5.392            // 1697
        ,   1.68    , -5.569            // 1698
        ,   1.68    , -5.392            // 1699
        ,  1.503    , -5.039            // 1700
        ,  1.503    , -5.216            // 1701
        ,   1.68    , -5.039            // 1702
        ,   1.68    , -5.216            // 1703
        ,  2.033    , -5.569            // 1704
        ,  2.033    , -5.392            // 1705
        ,  1.856    , -5.569            // 1706
        ,  1.856    , -5.392            // 1707
        ,  2.033    , -5.039            // 1708
        ,  2.033    , -5.216            // 1709
        ,  1.856    , -5.039            // 1710
        ,  1.856    , -5.216            // 1711
        ,  1.503    , -4.332            // 1712
        ,  1.503    , -4.508            // 1713
        ,   1.68    , -4.332            // 1714
        ,   1.68    , -4.508            // 1715
        ,  1.503    , -4.862            // 1716
        ,  1.503    , -4.685            // 1717
        ,   1.68    , -4.862            // 1718
        ,   1.68    , -4.685            // 1719
        ,  2.033    , -4.332            // 1720
        ,  2.033    , -4.508            // 1721
        ,  1.856    , -4.332            // 1722
        ,  1.856    , -4.508            // 1723
        ,  2.033    , -4.862            // 1724
        ,  2.033    , -4.685            // 1725
        ,  1.856    , -4.862            // 1726
        ,  1.856    , -4.685            // 1727
        ,   2.74    , -2.917            // 1728
        ,   2.74    , -3.094            // 1729
        ,  2.564    , -2.917            // 1730
        ,  2.564    , -3.094            // 1731
        ,   2.74    , -3.448            // 1732
        ,   2.74    , -3.271            // 1733
        ,  2.564    , -3.448            // 1734
        ,  2.564    , -3.271            // 1735
        ,   2.21    , -2.917            // 1736
        ,   2.21    , -3.094            // 1737
        ,  2.387    , -2.917            // 1738
        ,  2.387    , -3.094            // 1739
        ,   2.21    , -3.448            // 1740
        ,   2.21    , -3.271            // 1741
        ,  2.387    , -3.448            // 1742
        ,  2.387    , -3.271            // 1743
        ,   2.74    , -4.155            // 1744
        ,   2.74    , -3.978            // 1745
        ,  2.564    , -4.155            // 1746
        ,  2.564    , -3.978            // 1747
        ,   2.74    , -3.624            // 1748
        ,   2.74    , -3.801            // 1749
        ,  2.564    , -3.624            // 1750
        ,  2.564    , -3.801            // 1751
        ,   2.21    , -4.155            // 1752
        ,   2.21    , -3.978            // 1753
        ,  2.387    , -4.155            // 1754
        ,  2.387    , -3.978            // 1755
        ,   2.21    , -3.624            // 1756
        ,   2.21    , -3.801            // 1757
        ,  2.387    , -3.624            // 1758
        ,  2.387    , -3.801            // 1759
        ,  1.503    , -2.917            // 1760
        ,  1.503    , -3.094            // 1761
        ,   1.68    , -2.917            // 1762
        ,   1.68    , -3.094            // 1763
        ,  1.503    , -3.448            // 1764
        ,  1.503    , -3.271            // 1765
        ,   1.68    , -3.448            // 1766
        ,   1.68    , -3.271            // 1767
        ,  2.033    , -2.917            // 1768
        ,  2.033    , -3.094            // 1769
        ,  1.856    , -2.917            // 1770
        ,  1.856    , -3.094            // 1771
        ,  2.033    , -3.448            // 1772
        ,  2.033    , -3.271            // 1773
        ,  1.856    , -3.448            // 1774
        ,  1.856    , -3.271            // 1775
        ,  1.503    , -4.155            // 1776
        ,  1.503    , -3.978            // 1777
        ,   1.68    , -4.155            // 1778
        ,   1.68    , -3.978            // 1779
        ,  1.503    , -3.624            // 1780
        ,  1.503    , -3.801            // 1781
        ,   1.68    , -3.624            // 1782
        ,   1.68    , -3.801            // 1783
        ,  2.033    , -4.155            // 1784
        ,  2.033    , -3.978            // 1785
        ,  1.856    , -4.155            // 1786
        ,  1.856    , -3.978            // 1787
        ,  2.033    , -3.624            // 1788
        ,  2.033    , -3.801            // 1789
        ,  1.856    , -3.624            // 1790
        ,  1.856    , -3.801            // 1791
        ,  0.088    , -0.088            // 1792
        ,  0.088    , -0.265            // 1793
        ,  0.265    , -0.088            // 1794
        ,  0.265    , -0.265            // 1795
        ,  0.088    , -0.619            // 1796
        ,  0.088    , -0.442            // 1797
        ,  0.265    , -0.619            // 1798
        ,  0.265    , -0.442            // 1799
        ,  0.619    , -0.088            // 1800
        ,  0.619    , -0.265            // 1801
        ,  0.442    , -0.088            // 1802
        ,  0.442    , -0.265            // 1803
        ,  0.619    , -0.619            // 1804
        ,  0.619    , -0.442            // 1805
        ,  0.442    , -0.619            // 1806
        ,  0.442    , -0.442            // 1807
        ,  0.088    , -1.326            // 1808
        ,  0.088    , -1.149            // 1809
        ,  0.265    , -1.326            // 1810
        ,  0.265    , -1.149            // 1811
        ,  0.088    , -0.796            // 1812
        ,  0.088    , -0.972            // 1813
        ,  0.265    , -0.796            // 1814
        ,  0.265    , -0.972            // 1815
        ,  0.619    , -1.326            // 1816
        ,  0.619    , -1.149            // 1817
        ,  0.442    , -1.326            // 1818
        ,  0.442    , -1.149            // 1819
        ,  0.619    , -0.796            // 1820
        ,  0.619    , -0.972            // 1821
        ,  0.442    , -0.796            // 1822
        ,  0.442    , -0.972            // 1823
        ,  1.326    , -0.088            // 1824
        ,  1.326    , -0.265            // 1825
        ,  1.149    , -0.088            // 1826
        ,  1.149    , -0.265            // 1827
        ,  1.326    , -0.619            // 1828
        ,  1.326    , -0.442            // 1829
        ,  1.149    , -0.619            // 1830
        ,  1.149    , -0.442            // 1831
        ,  0.796    , -0.088            // 1832
        ,  0.796    , -0.265            // 1833
        ,  0.972    , -0.088            // 1834
        ,  0.972    , -0.265            // 1835
        ,  0.796    , -0.619            // 1836
        ,  0.796    , -0.442            // 1837
        ,  0.972    , -0.619            // 1838
        ,  0.972    , -0.442            // 1839
        ,  1.326    , -1.326            // 1840
        ,  1.326    , -1.149            // 1841
        ,  1.149    , -1.326            // 1842
        ,  1.149    , -1.149            // 1843
        ,  1.326    , -0.796            // 1844
        ,  1.326    , -0.972            // 1845
        ,  1.149    , -0.796            // 1846
        ,  1.149    , -0.972            // 1847
        ,  0.796    , -1.326            // 1848
        ,  0.796    , -1.149            // 1849
        ,  0.972    , -1.326            // 1850
        ,  0.972    , -1.149            // 1851
        ,  0.796    , -0.796            // 1852
        ,  0.796    , -0.972            // 1853
        ,  0.972    , -0.796            // 1854
        ,  0.972    , -0.972            // 1855
        ,  0.088    ,  -2.74            // 1856
        ,  0.088    , -2.564            // 1857
        ,  0.265    ,  -2.74            // 1858
        ,  0.265    , -2.564            // 1859
        ,  0.088    ,  -2.21            // 1860
        ,  0.088    , -2.387            // 1861
        ,  0.265    ,  -2.21            // 1862
        ,  0.265    , -2.387            // 1863
        ,  0.619    ,  -2.74            // 1864
        ,  0.619    , -2.564            // 1865
        ,  0.442    ,  -2.74            // 1866
        ,  0.442    , -2.564            // 1867
        ,  0.619    ,  -2.21            // 1868
        ,  0.619    , -2.387            // 1869
        ,  0.442    ,  -2.21            // 1870
        ,  0.442    , -2.387            // 1871
        ,  0.088    , -1.503            // 1872
        ,  0.088    ,  -1.68            // 1873
        ,  0.265    , -1.503            // 1874
        ,  0.265    ,  -1.68            // 1875
        ,  0.088    , -2.033            // 1876
        ,  0.088    , -1.856            // 1877
        ,  0.265    , -2.033            // 1878
        ,  0.265    , -1.856            // 1879
        ,  0.619    , -1.503            // 1880
        ,  0.619    ,  -1.68            // 1881
        ,  0.442    , -1.503            // 1882
        ,  0.442    ,  -1.68            // 1883
        ,  0.619    , -2.033            // 1884
        ,  0.619    , -1.856            // 1885
        ,  0.442    , -2.033            // 1886
        ,  0.442    , -1.856            // 1887
        ,  1.326    ,  -2.74            // 1888
        ,  1.326    , -2.564            // 1889
        ,  1.149    ,  -2.74            // 1890
        ,  1.149    , -2.564            // 1891
        ,  1.326    ,  -2.21            // 1892
        ,  1.326    , -2.387            // 1893
        ,  1.149    ,  -2.21            // 1894
        ,  1.149    , -2.387            // 1895
        ,  0.796    ,  -2.74            // 1896
        ,  0.796    , -2.564            // 1897
        ,  0.972    ,  -2.74            // 1898
        ,  0.972    , -2.564            // 1899
        ,  0.796    ,  -2.21            // 1900
        ,  0.796    , -2.387            // 1901
        ,  0.972    ,  -2.21            // 1902
        ,  0.972    , -2.387            // 1903
        ,  1.326    , -1.503            // 1904
        ,  1.326    ,  -1.68            // 1905
        ,  1.149    , -1.503            // 1906
        ,  1.149    ,  -1.68            // 1907
        ,  1.326    , -2.033            // 1908
        ,  1.326    , -1.856            // 1909
        ,  1.149    , -2.033            // 1910
        ,  1.149    , -1.856            // 1911
        ,  0.796    , -1.503            // 1912
        ,  0.796    ,  -1.68            // 1913
        ,  0.972    , -1.503            // 1914
        ,  0.972    ,  -1.68            // 1915
        ,  0.796    , -2.033            // 1916
        ,  0.796    , -1.856            // 1917
        ,  0.972    , -2.033            // 1918
        ,  0.972    , -1.856            // 1919
        ,   2.74    , -0.088            // 1920
        ,   2.74    , -0.265            // 1921
        ,  2.564    , -0.088            // 1922
        ,  2.564    , -0.265            // 1923
        ,   2.74    , -0.619            // 1924
        ,   2.74    , -0.442            // 1925
        ,  2.564    , -0.619            // 1926
        ,  2.564    , -0.442            // 1927
        ,   2.21    , -0.088            // 1928
        ,   2.21    , -0.265            // 1929
        ,  2.387    , -0.088            // 1930
        ,  2.387    , -0.265            // 1931
        ,   2.21    , -0.619            // 1932
        ,   2.21    , -0.442            // 1933
        ,  2.387    , -0.619            // 1934
        ,  2.387    , -0.442            // 1935
        ,   2.74    , -1.326            // 1936
        ,   2.74    , -1.149            // 1937
        ,  2.564    , -1.326            // 1938
        ,  2.564    , -1.149            // 1939
        ,   2.74    , -0.796            // 1940
        ,   2.74    , -0.972            // 1941
        ,  2.564    , -0.796            // 1942
        ,  2.564    , -0.972            // 1943
        ,   2.21    , -1.326            // 1944
        ,   2.21    , -1.149            // 1945
        ,  2.387    , -1.326            // 1946
        ,  2.387    , -1.149            // 1947
        ,   2.21    , -0.796            // 1948
        ,   2.21    , -0.972            // 1949
        ,  2.387    , -0.796            // 1950
        ,  2.387    , -0.972            // 1951
        ,  1.503    , -0.088            // 1952
        ,  1.503    , -0.265            // 1953
        ,   1.68    , -0.088            // 1954
        ,   1.68    , -0.265            // 1955
        ,  1.503    , -0.619            // 1956
        ,  1.503    , -0.442            // 1957
        ,   1.68    , -0.619            // 1958
        ,   1.68    , -0.442            // 1959
        ,  2.033    , -0.088            // 1960
        ,  2.033    , -0.265            // 1961
        ,  1.856    , -0.088            // 1962
        ,  1.856    , -0.265            // 1963
        ,  2.033    , -0.619            // 1964
        ,  2.033    , -0.442            // 1965
        ,  1.856    , -0.619            // 1966
        ,  1.856    , -0.442            // 1967
        ,  1.503    , -1.326            // 1968
        ,  1.503    , -1.149            // 1969
        ,   1.68    , -1.326            // 1970
        ,   1.68    , -1.149            // 1971
        ,  1.503    , -0.796            // 1972
        ,  1.503    , -0.972            // 1973
        ,   1.68    , -0.796            // 1974
        ,   1.68    , -0.972            // 1975
        ,  2.033    , -1.326            // 1976
        ,  2.033    , -1.149            // 1977
        ,  1.856    , -1.326            // 1978
        ,  1.856    , -1.149            // 1979
        ,  2.033    , -0.796            // 1980
        ,  2.033    , -0.972            // 1981
        ,  1.856    , -0.796            // 1982
        ,  1.856    , -0.972            // 1983
        ,   2.74    ,  -2.74            // 1984
        ,   2.74    , -2.564            // 1985
        ,  2.564    ,  -2.74            // 1986
        ,  2.564    , -2.564            // 1987
        ,   2.74    ,  -2.21            // 1988
        ,   2.74    , -2.387            // 1989
        ,  2.564    ,  -2.21            // 1990
        ,  2.564    , -2.387            // 1991
        ,   2.21    ,  -2.74            // 1992
        ,   2.21    , -2.564            // 1993
        ,  2.387    ,  -2.74            // 1994
        ,  2.387    , -2.564            // 1995
        ,   2.21    ,  -2.21            // 1996
        ,   2.21    , -2.387            // 1997
        ,  2.387    ,  -2.21            // 1998
        ,  2.387    , -2.387            // 1999
        ,   2.74    , -1.503            // 2000
        ,   2.74    ,  -1.68            // 2001
        ,  2.564    , -1.503            // 2002
        ,  2.564    ,  -1.68            // 2003
        ,   2.74    , -2.033            // 2004
        ,   2.74    , -1.856            // 2005
        ,  2.564    , -2.033            // 2006
        ,  2.564    , -1.856            // 2007
        ,   2.21    , -1.503            // 2008
        ,   2.21    ,  -1.68            // 2009
        ,  2.387    , -1.503            // 2010
        ,  2.387    ,  -1.68            // 2011
        ,   2.21    , -2.033            // 2012
        ,   2.21    , -1.856            // 2013
        ,  2.387    , -2.033            // 2014
        ,  2.387    , -1.856            // 2015
        ,  1.503    ,  -2.74            // 2016
        ,  1.503    , -2.564            // 2017
        ,   1.68    ,  -2.74            // 2018
        ,   1.68    , -2.564            // 2019
        ,  1.503    ,  -2.21            // 2020
        ,  1.503    , -2.387            // 2021
        ,   1.68    ,  -2.21            // 2022
        ,   1.68    , -2.387            // 2023
        ,  2.033    ,  -2.74            // 2024
        ,  2.033    , -2.564            // 2025
        ,  1.856    ,  -2.74            // 2026
        ,  1.856    , -2.564            // 2027
        ,  2.033    ,  -2.21            // 2028
        ,  2.033    , -2.387            // 2029
        ,  1.856    ,  -2.21            // 2030
        ,  1.856    , -2.387            // 2031
        ,  1.503    , -1.503            // 2032
        ,  1.503    ,  -1.68            // 2033
        ,   1.68    , -1.503            // 2034
        ,   1.68    ,  -1.68            // 2035
        ,  1.503    , -2.033            // 2036
        ,  1.503    , -1.856            // 2037
        ,   1.68    , -2.033            // 2038
        ,   1.68    , -1.856            // 2039
        ,  2.033    , -1.503            // 2040
        ,  2.033    ,  -1.68            // 2041
        ,  1.856    , -1.503            // 2042
        ,  1.856    ,  -1.68            // 2043
        ,  2.033    , -2.033            // 2044
        ,  2.033    , -1.856            // 2045
        ,  1.856    , -2.033            // 2046
        ,  1.856    , -1.856            // 2047
        , -5.569    ,  5.569            // 2048
        , -5.569    ,  5.392            // 2049
        , -5.392    ,  5.569            // 2050
        , -5.392    ,  5.392            // 2051
        , -5.569    ,  5.039            // 2052
        , -5.569    ,  5.216            // 2053
        , -5.392    ,  5.039            // 2054
        , -5.392    ,  5.216            // 2055
        , -5.039    ,  5.569            // 2056
        , -5.039    ,  5.392            // 2057
        , -5.216    ,  5.569            // 2058
        , -5.216    ,  5.392            // 2059
        , -5.039    ,  5.039            // 2060
        , -5.039    ,  5.216            // 2061
        , -5.216    ,  5.039            // 2062
        , -5.216    ,  5.216            // 2063
        , -5.569    ,  4.332            // 2064
        , -5.569    ,  4.508            // 2065
        , -5.392    ,  4.332            // 2066
        , -5.392    ,  4.508            // 2067
        , -5.569    ,  4.862            // 2068
        , -5.569    ,  4.685            // 2069
        , -5.392    ,  4.862            // 2070
        , -5.392    ,  4.685            // 2071
        , -5.039    ,  4.332            // 2072
        , -5.039    ,  4.508            // 2073
        , -5.216    ,  4.332            // 2074
        , -5.216    ,  4.508            // 2075
        , -5.039    ,  4.862            // 2076
        , -5.039    ,  4.685            // 2077
        , -5.216    ,  4.862            // 2078
        , -5.216    ,  4.685            // 2079
        , -4.332    ,  5.569            // 2080
        , -4.332    ,  5.392            // 2081
        , -4.508    ,  5.569            // 2082
        , -4.508    ,  5.392            // 2083
        , -4.332    ,  5.039            // 2084
        , -4.332    ,  5.216            // 2085
        , -4.508    ,  5.039            // 2086
        , -4.508    ,  5.216            // 2087
        , -4.862    ,  5.569            // 2088
        , -4.862    ,  5.392            // 2089
        , -4.685    ,  5.569            // 2090
        , -4.685    ,  5.392            // 2091
        , -4.862    ,  5.039            // 2092
        , -4.862    ,  5.216            // 2093
        , -4.685    ,  5.039            // 2094
        , -4.685    ,  5.216            // 2095
        , -4.332    ,  4.332            // 2096
        , -4.332    ,  4.508            // 2097
        , -4.508    ,  4.332            // 2098
        , -4.508    ,  4.508            // 2099
        , -4.332    ,  4.862            // 2100
        , -4.332    ,  4.685            // 2101
        , -4.508    ,  4.862            // 2102
        , -4.508    ,  4.685            // 2103
        , -4.862    ,  4.332            // 2104
        , -4.862    ,  4.508            // 2105
        , -4.685    ,  4.332            // 2106
        , -4.685    ,  4.508            // 2107
        , -4.862    ,  4.862            // 2108
        , -4.862    ,  4.685            // 2109
        , -4.685    ,  4.862            // 2110
        , -4.685    ,  4.685            // 2111
        , -5.569    ,  2.917            // 2112
        , -5.569    ,  3.094            // 2113
        , -5.392    ,  2.917            // 2114
        , -5.392    ,  3.094            // 2115
        , -5.569    ,  3.448            // 2116
        , -5.569    ,  3.271            // 2117
        , -5.392    ,  3.448            // 2118
        , -5.392    ,  3.271            // 2119
        , -5.039    ,  2.917            // 2120
        , -5.039    ,  3.094            // 2121
        , -5.216    ,  2.917            // 2122
        , -5.216    ,  3.094            // 2123
        , -5.039    ,  3.448            // 2124
        , -5.039    ,  3.271            // 2125
        , -5.216    ,  3.448            // 2126
        , -5.216    ,  3.271            // 2127
        , -5.569    ,  4.155            // 2128
        , -5.569    ,  3.978            // 2129
        , -5.392    ,  4.155            // 2130
        , -5.392    ,  3.978            // 2131
        , -5.569    ,  3.624            // 2132
        , -5.569    ,  3.801            // 2133
        , -5.392    ,  3.624            // 2134
        , -5.392    ,  3.801            // 2135
        , -5.039    ,  4.155            // 2136
        , -5.039    ,  3.978            // 2137
        , -5.216    ,  4.155            // 2138
        , -5.216    ,  3.978            // 2139
        , -5.039    ,  3.624            // 2140
        , -5.039    ,  3.801            // 2141
        , -5.216    ,  3.624            // 2142
        , -5.216    ,  3.801            // 2143
        , -4.332    ,  2.917            // 2144
        , -4.332    ,  3.094            // 2145
        , -4.508    ,  2.917            // 2146
        , -4.508    ,  3.094            // 2147
        , -4.332    ,  3.448            // 2148
        , -4.332    ,  3.271            // 2149
        , -4.508    ,  3.448            // 2150
        , -4.508    ,  3.271            // 2151
        , -4.862    ,  2.917            // 2152
        , -4.862    ,  3.094            // 2153
        , -4.685    ,  2.917            // 2154
        , -4.685    ,  3.094            // 2155
        , -4.862    ,  3.448            // 2156
        , -4.862    ,  3.271            // 2157
        , -4.685    ,  3.448            // 2158
        , -4.685    ,  3.271            // 2159
        , -4.332    ,  4.155            // 2160
        , -4.332    ,  3.978            // 2161
        , -4.508    ,  4.155            // 2162
        , -4.508    ,  3.978            // 2163
        , -4.332    ,  3.624            // 2164
        , -4.332    ,  3.801            // 2165
        , -4.508    ,  3.624            // 2166
        , -4.508    ,  3.801            // 2167
        , -4.862    ,  4.155            // 2168
        , -4.862    ,  3.978            // 2169
        , -4.685    ,  4.155            // 2170
        , -4.685    ,  3.978            // 2171
        , -4.862    ,  3.624            // 2172
        , -4.862    ,  3.801            // 2173
        , -4.685    ,  3.624            // 2174
        , -4.685    ,  3.801            // 2175
        , -2.917    ,  5.569            // 2176
        , -2.917    ,  5.392            // 2177
        , -3.094    ,  5.569            // 2178
        , -3.094    ,  5.392            // 2179
        , -2.917    ,  5.039            // 2180
        , -2.917    ,  5.216            // 2181
        , -3.094    ,  5.039            // 2182
        , -3.094    ,  5.216            // 2183
        , -3.448    ,  5.569            // 2184
        , -3.448    ,  5.392            // 2185
        , -3.271    ,  5.569            // 2186
        , -3.271    ,  5.392            // 2187
        , -3.448    ,  5.039            // 2188
        , -3.448    ,  5.216            // 2189
        , -3.271    ,  5.039            // 2190
        , -3.271    ,  5.216            // 2191
        , -2.917    ,  4.332            // 2192
        , -2.917    ,  4.508            // 2193
        , -3.094    ,  4.332            // 2194
        , -3.094    ,  4.508            // 2195
        , -2.917    ,  4.862            // 2196
        , -2.917    ,  4.685            // 2197
        , -3.094    ,  4.862            // 2198
        , -3.094    ,  4.685            // 2199
        , -3.448    ,  4.332            // 2200
        , -3.448    ,  4.508            // 2201
        , -3.271    ,  4.332            // 2202
        , -3.271    ,  4.508            // 2203
        , -3.448    ,  4.862            // 2204
        , -3.448    ,  4.685            // 2205
        , -3.271    ,  4.862            // 2206
        , -3.271    ,  4.685            // 2207
        , -4.155    ,  5.569            // 2208
        , -4.155    ,  5.392            // 2209
        , -3.978    ,  5.569            // 2210
        , -3.978    ,  5.392            // 2211
        , -4.155    ,  5.039            // 2212
        , -4.155    ,  5.216            // 2213
        , -3.978    ,  5.039            // 2214
        , -3.978    ,  5.216            // 2215
        , -3.624    ,  5.569            // 2216
        , -3.624    ,  5.392            // 2217
        , -3.801    ,  5.569            // 2218
        , -3.801    ,  5.392            // 2219
        , -3.624    ,  5.039            // 2220
        , -3.624    ,  5.216            // 2221
        , -3.801    ,  5.039            // 2222
        , -3.801    ,  5.216            // 2223
        , -4.155    ,  4.332            // 2224
        , -4.155    ,  4.508            // 2225
        , -3.978    ,  4.332            // 2226
        , -3.978    ,  4.508            // 2227
        , -4.155    ,  4.862            // 2228
        , -4.155    ,  4.685            // 2229
        , -3.978    ,  4.862            // 2230
        , -3.978    ,  4.685            // 2231
        , -3.624    ,  4.332            // 2232
        , -3.624    ,  4.508            // 2233
        , -3.801    ,  4.332            // 2234
        , -3.801    ,  4.508            // 2235
        , -3.624    ,  4.862            // 2236
        , -3.624    ,  4.685            // 2237
        , -3.801    ,  4.862            // 2238
        , -3.801    ,  4.685            // 2239
        , -2.917    ,  2.917            // 2240
        , -2.917    ,  3.094            // 2241
        , -3.094    ,  2.917            // 2242
        , -3.094    ,  3.094            // 2243
        , -2.917    ,  3.448            // 2244
        , -2.917    ,  3.271            // 2245
        , -3.094    ,  3.448            // 2246
        , -3.094    ,  3.271            // 2247
        , -3.448    ,  2.917            // 2248
        , -3.448    ,  3.094            // 2249
        , -3.271    ,  2.917            // 2250
        , -3.271    ,  3.094            // 2251
        , -3.448    ,  3.448            // 2252
        , -3.448    ,  3.271            // 2253
        , -3.271    ,  3.448            // 2254
        , -3.271    ,  3.271            // 2255
        , -2.917    ,  4.155            // 2256
        , -2.917    ,  3.978            // 2257
        , -3.094    ,  4.155            // 2258
        , -3.094    ,  3.978            // 2259
        , -2.917    ,  3.624            // 2260
        , -2.917    ,  3.801            // 2261
        , -3.094    ,  3.624            // 2262
        , -3.094    ,  3.801            // 2263
        , -3.448    ,  4.155            // 2264
        , -3.448    ,  3.978            // 2265
        , -3.271    ,  4.155            // 2266
        , -3.271    ,  3.978            // 2267
        , -3.448    ,  3.624            // 2268
        , -3.448    ,  3.801            // 2269
        , -3.271    ,  3.624            // 2270
        , -3.271    ,  3.801            // 2271
        , -4.155    ,  2.917            // 2272
        , -4.155    ,  3.094            // 2273
        , -3.978    ,  2.917            // 2274
        , -3.978    ,  3.094            // 2275
        , -4.155    ,  3.448            // 2276
        , -4.155    ,  3.271            // 2277
        , -3.978    ,  3.448            // 2278
        , -3.978    ,  3.271            // 2279
        , -3.624    ,  2.917            // 2280
        , -3.624    ,  3.094            // 2281
        , -3.801    ,  2.917            // 2282
        , -3.801    ,  3.094            // 2283
        , -3.624    ,  3.448            // 2284
        , -3.624    ,  3.271            // 2285
        , -3.801    ,  3.448            // 2286
        , -3.801    ,  3.271            // 2287
        , -4.155    ,  4.155            // 2288
        , -4.155    ,  3.978            // 2289
        , -3.978    ,  4.155            // 2290
        , -3.978    ,  3.978            // 2291
        , -4.155    ,  3.624            // 2292
        , -4.155    ,  3.801            // 2293
        , -3.978    ,  3.624            // 2294
        , -3.978    ,  3.801            // 2295
        , -3.624    ,  4.155            // 2296
        , -3.624    ,  3.978            // 2297
        , -3.801    ,  4.155            // 2298
        , -3.801    ,  3.978            // 2299
        , -3.624    ,  3.624            // 2300
        , -3.624    ,  3.801            // 2301
        , -3.801    ,  3.624            // 2302
        , -3.801    ,  3.801            // 2303
        , -5.569    ,  0.088            // 2304
        , -5.569    ,  0.265            // 2305
        , -5.392    ,  0.088            // 2306
        , -5.392    ,  0.265            // 2307
        , -5.569    ,  0.619            // 2308
        , -5.569    ,  0.442            // 2309
        , -5.392    ,  0.619            // 2310
        , -5.392    ,  0.442            // 2311
        , -5.039    ,  0.088            // 2312
        , -5.039    ,  0.265            // 2313
        , -5.216    ,  0.088            // 2314
        , -5.216    ,  0.265            // 2315
        , -5.039    ,  0.619            // 2316
        , -5.039    ,  0.442            // 2317
        , -5.216    ,  0.619            // 2318
        , -5.216    ,  0.442            // 2319
        , -5.569    ,  1.326            // 2320
        , -5.569    ,  1.149            // 2321
        , -5.392    ,  1.326            // 2322
        , -5.392    ,  1.149            // 2323
        , -5.569    ,  0.796            // 2324
        , -5.569    ,  0.972            // 2325
        , -5.392    ,  0.796            // 2326
        , -5.392    ,  0.972            // 2327
        , -5.039    ,  1.326            // 2328
        , -5.039    ,  1.149            // 2329
        , -5.216    ,  1.326            // 2330
        , -5.216    ,  1.149            // 2331
        , -5.039    ,  0.796            // 2332
        , -5.039    ,  0.972            // 2333
        , -5.216    ,  0.796            // 2334
        , -5.216    ,  0.972            // 2335
        , -4.332    ,  0.088            // 2336
        , -4.332    ,  0.265            // 2337
        , -4.508    ,  0.088            // 2338
        , -4.508    ,  0.265            // 2339
        , -4.332    ,  0.619            // 2340
        , -4.332    ,  0.442            // 2341
        , -4.508    ,  0.619            // 2342
        , -4.508    ,  0.442            // 2343
        , -4.862    ,  0.088            // 2344
        , -4.862    ,  0.265            // 2345
        , -4.685    ,  0.088            // 2346
        , -4.685    ,  0.265            // 2347
        , -4.862    ,  0.619            // 2348
        , -4.862    ,  0.442            // 2349
        , -4.685    ,  0.619            // 2350
        , -4.685    ,  0.442            // 2351
        , -4.332    ,  1.326            // 2352
        , -4.332    ,  1.149            // 2353
        , -4.508    ,  1.326            // 2354
        , -4.508    ,  1.149            // 2355
        , -4.332    ,  0.796            // 2356
        , -4.332    ,  0.972            // 2357
        , -4.508    ,  0.796            // 2358
        , -4.508    ,  0.972            // 2359
        , -4.862    ,  1.326            // 2360
        , -4.862    ,  1.149            // 2361
        , -4.685    ,  1.326            // 2362
        , -4.685    ,  1.149            // 2363
        , -4.862    ,  0.796            // 2364
        , -4.862    ,  0.972            // 2365
        , -4.685    ,  0.796            // 2366
        , -4.685    ,  0.972            // 2367
        , -5.569    ,   2.74            // 2368
        , -5.569    ,  2.564            // 2369
        , -5.392    ,   2.74            // 2370
        , -5.392    ,  2.564            // 2371
        , -5.569    ,   2.21            // 2372
        , -5.569    ,  2.387            // 2373
        , -5.392    ,   2.21            // 2374
        , -5.392    ,  2.387            // 2375
        , -5.039    ,   2.74            // 2376
        , -5.039    ,  2.564            // 2377
        , -5.216    ,   2.74            // 2378
        , -5.216    ,  2.564            // 2379
        , -5.039    ,   2.21            // 2380
        , -5.039    ,  2.387            // 2381
        , -5.216    ,   2.21            // 2382
        , -5.216    ,  2.387            // 2383
        , -5.569    ,  1.503            // 2384
        , -5.569    ,   1.68            // 2385
        , -5.392    ,  1.503            // 2386
        , -5.392    ,   1.68            // 2387
        , -5.569    ,  2.033            // 2388
        , -5.569    ,  1.856            // 2389
        , -5.392    ,  2.033            // 2390
        , -5.392    ,  1.856            // 2391
        , -5.039    ,  1.503            // 2392
        , -5.039    ,   1.68            // 2393
        , -5.216    ,  1.503            // 2394
        , -5.216    ,   1.68            // 2395
        , -5.039    ,  2.033            // 2396
        , -5.039    ,  1.856            // 2397
        , -5.216    ,  2.033            // 2398
        , -5.216    ,  1.856            // 2399
        , -4.332    ,   2.74            // 2400
        , -4.332    ,  2.564            // 2401
        , -4.508    ,   2.74            // 2402
        , -4.508    ,  2.564            // 2403
        , -4.332    ,   2.21            // 2404
        , -4.332    ,  2.387            // 2405
        , -4.508    ,   2.21            // 2406
        , -4.508    ,  2.387            // 2407
        , -4.862    ,   2.74            // 2408
        , -4.862    ,  2.564            // 2409
        , -4.685    ,   2.74            // 2410
        , -4.685    ,  2.564            // 2411
        , -4.862    ,   2.21            // 2412
        , -4.862    ,  2.387            // 2413
        , -4.685    ,   2.21            // 2414
        , -4.685    ,  2.387            // 2415
        , -4.332    ,  1.503            // 2416
        , -4.332    ,   1.68            // 2417
        , -4.508    ,  1.503            // 2418
        , -4.508    ,   1.68            // 2419
        , -4.332    ,  2.033            // 2420
        , -4.332    ,  1.856            // 2421
        , -4.508    ,  2.033            // 2422
        , -4.508    ,  1.856            // 2423
        , -4.862    ,  1.503            // 2424
        , -4.862    ,   1.68            // 2425
        , -4.685    ,  1.503            // 2426
        , -4.685    ,   1.68            // 2427
        , -4.862    ,  2.033            // 2428
        , -4.862    ,  1.856            // 2429
        , -4.685    ,  2.033            // 2430
        , -4.685    ,  1.856            // 2431
        , -2.917    ,  0.088            // 2432
        , -2.917    ,  0.265            // 2433
        , -3.094    ,  0.088            // 2434
        , -3.094    ,  0.265            // 2435
        , -2.917    ,  0.619            // 2436
        , -2.917    ,  0.442            // 2437
        , -3.094    ,  0.619            // 2438
        , -3.094    ,  0.442            // 2439
        , -3.448    ,  0.088            // 2440
        , -3.448    ,  0.265            // 2441
        , -3.271    ,  0.088            // 2442
        , -3.271    ,  0.265            // 2443
        , -3.448    ,  0.619            // 2444
        , -3.448    ,  0.442            // 2445
        , -3.271    ,  0.619            // 2446
        , -3.271    ,  0.442            // 2447
        , -2.917    ,  1.326            // 2448
        , -2.917    ,  1.149            // 2449
        , -3.094    ,  1.326            // 2450
        , -3.094    ,  1.149            // 2451
        , -2.917    ,  0.796            // 2452
        , -2.917    ,  0.972            // 2453
        , -3.094    ,  0.796            // 2454
        , -3.094    ,  0.972            // 2455
        , -3.448    ,  1.326            // 2456
        , -3.448    ,  1.149            // 2457
        , -3.271    ,  1.326            // 2458
        , -3.271    ,  1.149            // 2459
        , -3.448    ,  0.796            // 2460
        , -3.448    ,  0.972            // 2461
        , -3.271    ,  0.796            // 2462
        , -3.271    ,  0.972            // 2463
        , -4.155    ,  0.088            // 2464
        , -4.155    ,  0.265            // 2465
        , -3.978    ,  0.088            // 2466
        , -3.978    ,  0.265            // 2467
        , -4.155    ,  0.619            // 2468
        , -4.155    ,  0.442            // 2469
        , -3.978    ,  0.619            // 2470
        , -3.978    ,  0.442            // 2471
        , -3.624    ,  0.088            // 2472
        , -3.624    ,  0.265            // 2473
        , -3.801    ,  0.088            // 2474
        , -3.801    ,  0.265            // 2475
        , -3.624    ,  0.619            // 2476
        , -3.624    ,  0.442            // 2477
        , -3.801    ,  0.619            // 2478
        , -3.801    ,  0.442            // 2479
        , -4.155    ,  1.326            // 2480
        , -4.155    ,  1.149            // 2481
        , -3.978    ,  1.326            // 2482
        , -3.978    ,  1.149            // 2483
        , -4.155    ,  0.796            // 2484
        , -4.155    ,  0.972            // 2485
        , -3.978    ,  0.796            // 2486
        , -3.978    ,  0.972            // 2487
        , -3.624    ,  1.326            // 2488
        , -3.624    ,  1.149            // 2489
        , -3.801    ,  1.326            // 2490
        , -3.801    ,  1.149            // 2491
        , -3.624    ,  0.796            // 2492
        , -3.624    ,  0.972            // 2493
        , -3.801    ,  0.796            // 2494
        , -3.801    ,  0.972            // 2495
        , -2.917    ,   2.74            // 2496
        , -2.917    ,  2.564            // 2497
        , -3.094    ,   2.74            // 2498
        , -3.094    ,  2.564            // 2499
        , -2.917    ,   2.21            // 2500
        , -2.917    ,  2.387            // 2501
        , -3.094    ,   2.21            // 2502
        , -3.094    ,  2.387            // 2503
        , -3.448    ,   2.74            // 2504
        , -3.448    ,  2.564            // 2505
        , -3.271    ,   2.74            // 2506
        , -3.271    ,  2.564            // 2507
        , -3.448    ,   2.21            // 2508
        , -3.448    ,  2.387            // 2509
        , -3.271    ,   2.21            // 2510
        , -3.271    ,  2.387            // 2511
        , -2.917    ,  1.503            // 2512
        , -2.917    ,   1.68            // 2513
        , -3.094    ,  1.503            // 2514
        , -3.094    ,   1.68            // 2515
        , -2.917    ,  2.033            // 2516
        , -2.917    ,  1.856            // 2517
        , -3.094    ,  2.033            // 2518
        , -3.094    ,  1.856            // 2519
        , -3.448    ,  1.503            // 2520
        , -3.448    ,   1.68            // 2521
        , -3.271    ,  1.503            // 2522
        , -3.271    ,   1.68            // 2523
        , -3.448    ,  2.033            // 2524
        , -3.448    ,  1.856            // 2525
        , -3.271    ,  2.033            // 2526
        , -3.271    ,  1.856            // 2527
        , -4.155    ,   2.74            // 2528
        , -4.155    ,  2.564            // 2529
        , -3.978    ,   2.74            // 2530
        , -3.978    ,  2.564            // 2531
        , -4.155    ,   2.21            // 2532
        , -4.155    ,  2.387            // 2533
        , -3.978    ,   2.21            // 2534
        , -3.978    ,  2.387            // 2535
        , -3.624    ,   2.74            // 2536
        , -3.624    ,  2.564            // 2537
        , -3.801    ,   2.74            // 2538
        , -3.801    ,  2.564            // 2539
        , -3.624    ,   2.21            // 2540
        , -3.624    ,  2.387            // 2541
        , -3.801    ,   2.21            // 2542
        , -3.801    ,  2.387            // 2543
        , -4.155    ,  1.503            // 2544
        , -4.155    ,   1.68            // 2545
        , -3.978    ,  1.503            // 2546
        , -3.978    ,   1.68            // 2547
        , -4.155    ,  2.033            // 2548
        , -4.155    ,  1.856            // 2549
        , -3.978    ,  2.033            // 2550
        , -3.978    ,  1.856            // 2551
        , -3.624    ,  1.503            // 2552
        , -3.624    ,   1.68            // 2553
        , -3.801    ,  1.503            // 2554
        , -3.801    ,   1.68            // 2555
        , -3.624    ,  2.033            // 2556
        , -3.624    ,  1.856            // 2557
        , -3.801    ,  2.033            // 2558
        , -3.801    ,  1.856            // 2559
        , -0.088    ,  5.569            // 2560
        , -0.088    ,  5.392            // 2561
        , -0.265    ,  5.569            // 2562
        , -0.265    ,  5.392            // 2563
        , -0.088    ,  5.039            // 2564
        , -0.088    ,  5.216            // 2565
        , -0.265    ,  5.039            // 2566
        , -0.265    ,  5.216            // 2567
        , -0.619    ,  5.569            // 2568
        , -0.619    ,  5.392            // 2569
        , -0.442    ,  5.569            // 2570
        , -0.442    ,  5.392            // 2571
        , -0.619    ,  5.039            // 2572
        , -0.619    ,  5.216            // 2573
        , -0.442    ,  5.039            // 2574
        , -0.442    ,  5.216            // 2575
        , -0.088    ,  4.332            // 2576
        , -0.088    ,  4.508            // 2577
        , -0.265    ,  4.332            // 2578
        , -0.265    ,  4.508            // 2579
        , -0.088    ,  4.862            // 2580
        , -0.088    ,  4.685            // 2581
        , -0.265    ,  4.862            // 2582
        , -0.265    ,  4.685            // 2583
        , -0.619    ,  4.332            // 2584
        , -0.619    ,  4.508            // 2585
        , -0.442    ,  4.332            // 2586
        , -0.442    ,  4.508            // 2587
        , -0.619    ,  4.862            // 2588
        , -0.619    ,  4.685            // 2589
        , -0.442    ,  4.862            // 2590
        , -0.442    ,  4.685            // 2591
        , -1.326    ,  5.569            // 2592
        , -1.326    ,  5.392            // 2593
        , -1.149    ,  5.569            // 2594
        , -1.149    ,  5.392            // 2595
        , -1.326    ,  5.039            // 2596
        , -1.326    ,  5.216            // 2597
        , -1.149    ,  5.039            // 2598
        , -1.149    ,  5.216            // 2599
        , -0.796    ,  5.569            // 2600
        , -0.796    ,  5.392            // 2601
        , -0.972    ,  5.569            // 2602
        , -0.972    ,  5.392            // 2603
        , -0.796    ,  5.039            // 2604
        , -0.796    ,  5.216            // 2605
        , -0.972    ,  5.039            // 2606
        , -0.972    ,  5.216            // 2607
        , -1.326    ,  4.332            // 2608
        , -1.326    ,  4.508            // 2609
        , -1.149    ,  4.332            // 2610
        , -1.149    ,  4.508            // 2611
        , -1.326    ,  4.862            // 2612
        , -1.326    ,  4.685            // 2613
        , -1.149    ,  4.862            // 2614
        , -1.149    ,  4.685            // 2615
        , -0.796    ,  4.332            // 2616
        , -0.796    ,  4.508            // 2617
        , -0.972    ,  4.332            // 2618
        , -0.972    ,  4.508            // 2619
        , -0.796    ,  4.862            // 2620
        , -0.796    ,  4.685            // 2621
        , -0.972    ,  4.862            // 2622
        , -0.972    ,  4.685            // 2623
        , -0.088    ,  2.917            // 2624
        , -0.088    ,  3.094            // 2625
        , -0.265    ,  2.917            // 2626
        , -0.265    ,  3.094            // 2627
        , -0.088    ,  3.448            // 2628
        , -0.088    ,  3.271            // 2629
        , -0.265    ,  3.448            // 2630
        , -0.265    ,  3.271            // 2631
        , -0.619    ,  2.917            // 2632
        , -0.619    ,  3.094            // 2633
        , -0.442    ,  2.917            // 2634
        , -0.442    ,  3.094            // 2635
        , -0.619    ,  3.448            // 2636
        , -0.619    ,  3.271            // 2637
        , -0.442    ,  3.448            // 2638
        , -0.442    ,  3.271            // 2639
        , -0.088    ,  4.155            // 2640
        , -0.088    ,  3.978            // 2641
        , -0.265    ,  4.155            // 2642
        , -0.265    ,  3.978            // 2643
        , -0.088    ,  3.624            // 2644
        , -0.088    ,  3.801            // 2645
        , -0.265    ,  3.624            // 2646
        , -0.265    ,  3.801            // 2647
        , -0.619    ,  4.155            // 2648
        , -0.619    ,  3.978            // 2649
        , -0.442    ,  4.155            // 2650
        , -0.442    ,  3.978            // 2651
        , -0.619    ,  3.624            // 2652
        , -0.619    ,  3.801            // 2653
        , -0.442    ,  3.624            // 2654
        , -0.442    ,  3.801            // 2655
        , -1.326    ,  2.917            // 2656
        , -1.326    ,  3.094            // 2657
        , -1.149    ,  2.917            // 2658
        , -1.149    ,  3.094            // 2659
        , -1.326    ,  3.448            // 2660
        , -1.326    ,  3.271            // 2661
        , -1.149    ,  3.448            // 2662
        , -1.149    ,  3.271            // 2663
        , -0.796    ,  2.917            // 2664
        , -0.796    ,  3.094            // 2665
        , -0.972    ,  2.917            // 2666
        , -0.972    ,  3.094            // 2667
        , -0.796    ,  3.448            // 2668
        , -0.796    ,  3.271            // 2669
        , -0.972    ,  3.448            // 2670
        , -0.972    ,  3.271            // 2671
        , -1.326    ,  4.155            // 2672
        , -1.326    ,  3.978            // 2673
        , -1.149    ,  4.155            // 2674
        , -1.149    ,  3.978            // 2675
        , -1.326    ,  3.624            // 2676
        , -1.326    ,  3.801            // 2677
        , -1.149    ,  3.624            // 2678
        , -1.149    ,  3.801            // 2679
        , -0.796    ,  4.155            // 2680
        , -0.796    ,  3.978            // 2681
        , -0.972    ,  4.155            // 2682
        , -0.972    ,  3.978            // 2683
        , -0.796    ,  3.624            // 2684
        , -0.796    ,  3.801            // 2685
        , -0.972    ,  3.624            // 2686
        , -0.972    ,  3.801            // 2687
        ,  -2.74    ,  5.569            // 2688
        ,  -2.74    ,  5.392            // 2689
        , -2.564    ,  5.569            // 2690
        , -2.564    ,  5.392            // 2691
        ,  -2.74    ,  5.039            // 2692
        ,  -2.74    ,  5.216            // 2693
        , -2.564    ,  5.039            // 2694
        , -2.564    ,  5.216            // 2695
        ,  -2.21    ,  5.569            // 2696
        ,  -2.21    ,  5.392            // 2697
        , -2.387    ,  5.569            // 2698
        , -2.387    ,  5.392            // 2699
        ,  -2.21    ,  5.039            // 2700
        ,  -2.21    ,  5.216            // 2701
        , -2.387    ,  5.039            // 2702
        , -2.387    ,  5.216            // 2703
        ,  -2.74    ,  4.332            // 2704
        ,  -2.74    ,  4.508            // 2705
        , -2.564    ,  4.332            // 2706
        , -2.564    ,  4.508            // 2707
        ,  -2.74    ,  4.862            // 2708
        ,  -2.74    ,  4.685            // 2709
        , -2.564    ,  4.862            // 2710
        , -2.564    ,  4.685            // 2711
        ,  -2.21    ,  4.332            // 2712
        ,  -2.21    ,  4.508            // 2713
        , -2.387    ,  4.332            // 2714
        , -2.387    ,  4.508            // 2715
        ,  -2.21    ,  4.862            // 2716
        ,  -2.21    ,  4.685            // 2717
        , -2.387    ,  4.862            // 2718
        , -2.387    ,  4.685            // 2719
        , -1.503    ,  5.569            // 2720
        , -1.503    ,  5.392            // 2721
        ,  -1.68    ,  5.569            // 2722
        ,  -1.68    ,  5.392            // 2723
        , -1.503    ,  5.039            // 2724
        , -1.503    ,  5.216            // 2725
        ,  -1.68    ,  5.039            // 2726
        ,  -1.68    ,  5.216            // 2727
        , -2.033    ,  5.569            // 2728
        , -2.033    ,  5.392            // 2729
        , -1.856    ,  5.569            // 2730
        , -1.856    ,  5.392            // 2731
        , -2.033    ,  5.039            // 2732
        , -2.033    ,  5.216            // 2733
        , -1.856    ,  5.039            // 2734
        , -1.856    ,  5.216            // 2735
        , -1.503    ,  4.332            // 2736
        , -1.503    ,  4.508            // 2737
        ,  -1.68    ,  4.332            // 2738
        ,  -1.68    ,  4.508            // 2739
        , -1.503    ,  4.862            // 2740
        , -1.503    ,  4.685            // 2741
        ,  -1.68    ,  4.862            // 2742
        ,  -1.68    ,  4.685            // 2743
        , -2.033    ,  4.332            // 2744
        , -2.033    ,  4.508            // 2745
        , -1.856    ,  4.332            // 2746
        , -1.856    ,  4.508            // 2747
        , -2.033    ,  4.862            // 2748
        , -2.033    ,  4.685            // 2749
        , -1.856    ,  4.862            // 2750
        , -1.856    ,  4.685            // 2751
        ,  -2.74    ,  2.917            // 2752
        ,  -2.74    ,  3.094            // 2753
        , -2.564    ,  2.917            // 2754
        , -2.564    ,  3.094            // 2755
        ,  -2.74    ,  3.448            // 2756
        ,  -2.74    ,  3.271            // 2757
        , -2.564    ,  3.448            // 2758
        , -2.564    ,  3.271            // 2759
        ,  -2.21    ,  2.917            // 2760
        ,  -2.21    ,  3.094            // 2761
        , -2.387    ,  2.917            // 2762
        , -2.387    ,  3.094            // 2763
        ,  -2.21    ,  3.448            // 2764
        ,  -2.21    ,  3.271            // 2765
        , -2.387    ,  3.448            // 2766
        , -2.387    ,  3.271            // 2767
        ,  -2.74    ,  4.155            // 2768
        ,  -2.74    ,  3.978            // 2769
        , -2.564    ,  4.155            // 2770
        , -2.564    ,  3.978            // 2771
        ,  -2.74    ,  3.624            // 2772
        ,  -2.74    ,  3.801            // 2773
        , -2.564    ,  3.624            // 2774
        , -2.564    ,  3.801            // 2775
        ,  -2.21    ,  4.155            // 2776
        ,  -2.21    ,  3.978            // 2777
        , -2.387    ,  4.155            // 2778
        , -2.387    ,  3.978            // 2779
        ,  -2.21    ,  3.624            // 2780
        ,  -2.21    ,  3.801            // 2781
        , -2.387    ,  3.624            // 2782
        , -2.387    ,  3.801            // 2783
        , -1.503    ,  2.917            // 2784
        , -1.503    ,  3.094            // 2785
        ,  -1.68    ,  2.917            // 2786
        ,  -1.68    ,  3.094            // 2787
        , -1.503    ,  3.448            // 2788
        , -1.503    ,  3.271            // 2789
        ,  -1.68    ,  3.448            // 2790
        ,  -1.68    ,  3.271            // 2791
        , -2.033    ,  2.917            // 2792
        , -2.033    ,  3.094            // 2793
        , -1.856    ,  2.917            // 2794
        , -1.856    ,  3.094            // 2795
        , -2.033    ,  3.448            // 2796
        , -2.033    ,  3.271            // 2797
        , -1.856    ,  3.448            // 2798
        , -1.856    ,  3.271            // 2799
        , -1.503    ,  4.155            // 2800
        , -1.503    ,  3.978            // 2801
        ,  -1.68    ,  4.155            // 2802
        ,  -1.68    ,  3.978            // 2803
        , -1.503    ,  3.624            // 2804
        , -1.503    ,  3.801            // 2805
        ,  -1.68    ,  3.624            // 2806
        ,  -1.68    ,  3.801            // 2807
        , -2.033    ,  4.155            // 2808
        , -2.033    ,  3.978            // 2809
        , -1.856    ,  4.155            // 2810
        , -1.856    ,  3.978            // 2811
        , -2.033    ,  3.624            // 2812
        , -2.033    ,  3.801            // 2813
        , -1.856    ,  3.624            // 2814
        , -1.856    ,  3.801            // 2815
        , -0.088    ,  0.088            // 2816
        , -0.088    ,  0.265            // 2817
        , -0.265    ,  0.088            // 2818
        , -0.265    ,  0.265            // 2819
        , -0.088    ,  0.619            // 2820
        , -0.088    ,  0.442            // 2821
        , -0.265    ,  0.619            // 2822
        , -0.265    ,  0.442            // 2823
        , -0.619    ,  0.088            // 2824
        , -0.619    ,  0.265            // 2825
        , -0.442    ,  0.088            // 2826
        , -0.442    ,  0.265            // 2827
        , -0.619    ,  0.619            // 2828
        , -0.619    ,  0.442            // 2829
        , -0.442    ,  0.619            // 2830
        , -0.442    ,  0.442            // 2831
        , -0.088    ,  1.326            // 2832
        , -0.088    ,  1.149            // 2833
        , -0.265    ,  1.326            // 2834
        , -0.265    ,  1.149            // 2835
        , -0.088    ,  0.796            // 2836
        , -0.088    ,  0.972            // 2837
        , -0.265    ,  0.796            // 2838
        , -0.265    ,  0.972            // 2839
        , -0.619    ,  1.326            // 2840
        , -0.619    ,  1.149            // 2841
        , -0.442    ,  1.326            // 2842
        , -0.442    ,  1.149            // 2843
        , -0.619    ,  0.796            // 2844
        , -0.619    ,  0.972            // 2845
        , -0.442    ,  0.796            // 2846
        , -0.442    ,  0.972            // 2847
        , -1.326    ,  0.088            // 2848
        , -1.326    ,  0.265            // 2849
        , -1.149    ,  0.088            // 2850
        , -1.149    ,  0.265            // 2851
        , -1.326    ,  0.619            // 2852
        , -1.326    ,  0.442            // 2853
        , -1.149    ,  0.619            // 2854
        , -1.149    ,  0.442            // 2855
        , -0.796    ,  0.088            // 2856
        , -0.796    ,  0.265            // 2857
        , -0.972    ,  0.088            // 2858
        , -0.972    ,  0.265            // 2859
        , -0.796    ,  0.619            // 2860
        , -0.796    ,  0.442            // 2861
        , -0.972    ,  0.619            // 2862
        , -0.972    ,  0.442            // 2863
        , -1.326    ,  1.326            // 2864
        , -1.326    ,  1.149            // 2865
        , -1.149    ,  1.326            // 2866
        , -1.149    ,  1.149            // 2867
        , -1.326    ,  0.796            // 2868
        , -1.326    ,  0.972            // 2869
        , -1.149    ,  0.796            // 2870
        , -1.149    ,  0.972            // 2871
        , -0.796    ,  1.326            // 2872
        , -0.796    ,  1.149            // 2873
        , -0.972    ,  1.326            // 2874
        , -0.972    ,  1.149            // 2875
        , -0.796    ,  0.796            // 2876
        , -0.796    ,  0.972            // 2877
        , -0.972    ,  0.796            // 2878
        , -0.972    ,  0.972            // 2879
        , -0.088    ,   2.74            // 2880
        , -0.088    ,  2.564            // 2881
        , -0.265    ,   2.74            // 2882
        , -0.265    ,  2.564            // 2883
        , -0.088    ,   2.21            // 2884
        , -0.088    ,  2.387            // 2885
        , -0.265    ,   2.21            // 2886
        , -0.265    ,  2.387            // 2887
        , -0.619    ,   2.74            // 2888
        , -0.619    ,  2.564            // 2889
        , -0.442    ,   2.74            // 2890
        , -0.442    ,  2.564            // 2891
        , -0.619    ,   2.21            // 2892
        , -0.619    ,  2.387            // 2893
        , -0.442    ,   2.21            // 2894
        , -0.442    ,  2.387            // 2895
        , -0.088    ,  1.503            // 2896
        , -0.088    ,   1.68            // 2897
        , -0.265    ,  1.503            // 2898
        , -0.265    ,   1.68            // 2899
        , -0.088    ,  2.033            // 2900
        , -0.088    ,  1.856            // 2901
        , -0.265    ,  2.033            // 2902
        , -0.265    ,  1.856            // 2903
        , -0.619    ,  1.503            // 2904
        , -0.619    ,   1.68            // 2905
        , -0.442    ,  1.503            // 2906
        , -0.442    ,   1.68            // 2907
        , -0.619    ,  2.033            // 2908
        , -0.619    ,  1.856            // 2909
        , -0.442    ,  2.033            // 2910
        , -0.442    ,  1.856            // 2911
        , -1.326    ,   2.74            // 2912
        , -1.326    ,  2.564            // 2913
        , -1.149    ,   2.74            // 2914
        , -1.149    ,  2.564            // 2915
        , -1.326    ,   2.21            // 2916
        , -1.326    ,  2.387            // 2917
        , -1.149    ,   2.21            // 2918
        , -1.149    ,  2.387            // 2919
        , -0.796    ,   2.74            // 2920
        , -0.796    ,  2.564            // 2921
        , -0.972    ,   2.74            // 2922
        , -0.972    ,  2.564            // 2923
        , -0.796    ,   2.21            // 2924
        , -0.796    ,  2.387            // 2925
        , -0.972    ,   2.21            // 2926
        , -0.972    ,  2.387            // 2927
        , -1.326    ,  1.503            // 2928
        , -1.326    ,   1.68            // 2929
        , -1.149    ,  1.503            // 2930
        , -1.149    ,   1.68            // 2931
        , -1.326    ,  2.033            // 2932
        , -1.326    ,  1.856            // 2933
        , -1.149    ,  2.033            // 2934
        , -1.149    ,  1.856            // 2935
        , -0.796    ,  1.503            // 2936
        , -0.796    ,   1.68            // 2937
        , -0.972    ,  1.503            // 2938
        , -0.972    ,   1.68            // 2939
        , -0.796    ,  2.033            // 2940
        , -0.796    ,  1.856            // 2941
        , -0.972    ,  2.033            // 2942
        , -0.972    ,  1.856            // 2943
        ,  -2.74    ,  0.088            // 2944
        ,  -2.74    ,  0.265            // 2945
        , -2.564    ,  0.088            // 2946
        , -2.564    ,  0.265            // 2947
        ,  -2.74    ,  0.619            // 2948
        ,  -2.74    ,  0.442            // 2949
        , -2.564    ,  0.619            // 2950
        , -2.564    ,  0.442            // 2951
        ,  -2.21    ,  0.088            // 2952
        ,  -2.21    ,  0.265            // 2953
        , -2.387    ,  0.088            // 2954
        , -2.387    ,  0.265            // 2955
        ,  -2.21    ,  0.619            // 2956
        ,  -2.21    ,  0.442            // 2957
        , -2.387    ,  0.619            // 2958
        , -2.387    ,  0.442            // 2959
        ,  -2.74    ,  1.326            // 2960
        ,  -2.74    ,  1.149            // 2961
        , -2.564    ,  1.326            // 2962
        , -2.564    ,  1.149            // 2963
        ,  -2.74    ,  0.796            // 2964
        ,  -2.74    ,  0.972            // 2965
        , -2.564    ,  0.796            // 2966
        , -2.564    ,  0.972            // 2967
        ,  -2.21    ,  1.326            // 2968
        ,  -2.21    ,  1.149            // 2969
        , -2.387    ,  1.326            // 2970
        , -2.387    ,  1.149            // 2971
        ,  -2.21    ,  0.796            // 2972
        ,  -2.21    ,  0.972            // 2973
        , -2.387    ,  0.796            // 2974
        , -2.387    ,  0.972            // 2975
        , -1.503    ,  0.088            // 2976
        , -1.503    ,  0.265            // 2977
        ,  -1.68    ,  0.088            // 2978
        ,  -1.68    ,  0.265            // 2979
        , -1.503    ,  0.619            // 2980
        , -1.503    ,  0.442            // 2981
        ,  -1.68    ,  0.619            // 2982
        ,  -1.68    ,  0.442            // 2983
        , -2.033    ,  0.088            // 2984
        , -2.033    ,  0.265            // 2985
        , -1.856    ,  0.088            // 2986
        , -1.856    ,  0.265            // 2987
        , -2.033    ,  0.619            // 2988
        , -2.033    ,  0.442            // 2989
        , -1.856    ,  0.619            // 2990
        , -1.856    ,  0.442            // 2991
        , -1.503    ,  1.326            // 2992
        , -1.503    ,  1.149            // 2993
        ,  -1.68    ,  1.326            // 2994
        ,  -1.68    ,  1.149            // 2995
        , -1.503    ,  0.796            // 2996
        , -1.503    ,  0.972            // 2997
        ,  -1.68    ,  0.796            // 2998
        ,  -1.68    ,  0.972            // 2999
        , -2.033    ,  1.326            // 3000
        , -2.033    ,  1.149            // 3001
        , -1.856    ,  1.326            // 3002
        , -1.856    ,  1.149            // 3003
        , -2.033    ,  0.796            // 3004
        , -2.033    ,  0.972            // 3005
        , -1.856    ,  0.796            // 3006
        , -1.856    ,  0.972            // 3007
        ,  -2.74    ,   2.74            // 3008
        ,  -2.74    ,  2.564            // 3009
        , -2.564    ,   2.74            // 3010
        , -2.564    ,  2.564            // 3011
        ,  -2.74    ,   2.21            // 3012
        ,  -2.74    ,  2.387            // 3013
        , -2.564    ,   2.21            // 3014
        , -2.564    ,  2.387            // 3015
        ,  -2.21    ,   2.74            // 3016
        ,  -2.21    ,  2.564            // 3017
        , -2.387    ,   2.74            // 3018
        , -2.387    ,  2.564            // 3019
        ,  -2.21    ,   2.21            // 3020
        ,  -2.21    ,  2.387            // 3021
        , -2.387    ,   2.21            // 3022
        , -2.387    ,  2.387            // 3023
        ,  -2.74    ,  1.503            // 3024
        ,  -2.74    ,   1.68            // 3025
        , -2.564    ,  1.503            // 3026
        , -2.564    ,   1.68            // 3027
        ,  -2.74    ,  2.033            // 3028
        ,  -2.74    ,  1.856            // 3029
        , -2.564    ,  2.033            // 3030
        , -2.564    ,  1.856            // 3031
        ,  -2.21    ,  1.503            // 3032
        ,  -2.21    ,   1.68            // 3033
        , -2.387    ,  1.503            // 3034
        , -2.387    ,   1.68            // 3035
        ,  -2.21    ,  2.033            // 3036
        ,  -2.21    ,  1.856            // 3037
        , -2.387    ,  2.033            // 3038
        , -2.387    ,  1.856            // 3039
        , -1.503    ,   2.74            // 3040
        , -1.503    ,  2.564            // 3041
        ,  -1.68    ,   2.74            // 3042
        ,  -1.68    ,  2.564            // 3043
        , -1.503    ,   2.21            // 3044
        , -1.503    ,  2.387            // 3045
        ,  -1.68    ,   2.21            // 3046
        ,  -1.68    ,  2.387            // 3047
        , -2.033    ,   2.74            // 3048
        , -2.033    ,  2.564            // 3049
        , -1.856    ,   2.74            // 3050
        , -1.856    ,  2.564            // 3051
        , -2.033    ,   2.21            // 3052
        , -2.033    ,  2.387            // 3053
        , -1.856    ,   2.21            // 3054
        , -1.856    ,  2.387            // 3055
        , -1.503    ,  1.503            // 3056
        , -1.503    ,   1.68            // 3057
        ,  -1.68    ,  1.503            // 3058
        ,  -1.68    ,   1.68            // 3059
        , -1.503    ,  2.033            // 3060
        , -1.503    ,  1.856            // 3061
        ,  -1.68    ,  2.033            // 3062
        ,  -1.68    ,  1.856            // 3063
        , -2.033    ,  1.503            // 3064
        , -2.033    ,   1.68            // 3065
        , -1.856    ,  1.503            // 3066
        , -1.856    ,   1.68            // 3067
        , -2.033    ,  2.033            // 3068
        , -2.033    ,  1.856            // 3069
        , -1.856    ,  2.033            // 3070
        , -1.856    ,  1.856            // 3071
        , -5.569    , -5.569            // 3072
        , -5.569    , -5.392            // 3073
        , -5.392    , -5.569            // 3074
        , -5.392    , -5.392            // 3075
        , -5.569    , -5.039            // 3076
        , -5.569    , -5.216            // 3077
        , -5.392    , -5.039            // 3078
        , -5.392    , -5.216            // 3079
        , -5.039    , -5.569            // 3080
        , -5.039    , -5.392            // 3081
        , -5.216    , -5.569            // 3082
        , -5.216    , -5.392            // 3083
        , -5.039    , -5.039            // 3084
        , -5.039    , -5.216            // 3085
        , -5.216    , -5.039            // 3086
        , -5.216    , -5.216            // 3087
        , -5.569    , -4.332            // 3088
        , -5.569    , -4.508            // 3089
        , -5.392    , -4.332            // 3090
        , -5.392    , -4.508            // 3091
        , -5.569    , -4.862            // 3092
        , -5.569    , -4.685            // 3093
        , -5.392    , -4.862            // 3094
        , -5.392    , -4.685            // 3095
        , -5.039    , -4.332            // 3096
        , -5.039    , -4.508            // 3097
        , -5.216    , -4.332            // 3098
        , -5.216    , -4.508            // 3099
        , -5.039    , -4.862            // 3100
        , -5.039    , -4.685            // 3101
        , -5.216    , -4.862            // 3102
        , -5.216    , -4.685            // 3103
        , -4.332    , -5.569            // 3104
        , -4.332    , -5.392            // 3105
        , -4.508    , -5.569            // 3106
        , -4.508    , -5.392            // 3107
        , -4.332    , -5.039            // 3108
        , -4.332    , -5.216            // 3109
        , -4.508    , -5.039            // 3110
        , -4.508    , -5.216            // 3111
        , -4.862    , -5.569            // 3112
        , -4.862    , -5.392            // 3113
        , -4.685    , -5.569            // 3114
        , -4.685    , -5.392            // 3115
        , -4.862    , -5.039            // 3116
        , -4.862    , -5.216            // 3117
        , -4.685    , -5.039            // 3118
        , -4.685    , -5.216            // 3119
        , -4.332    , -4.332            // 3120
        , -4.332    , -4.508            // 3121
        , -4.508    , -4.332            // 3122
        , -4.508    , -4.508            // 3123
        , -4.332    , -4.862            // 3124
        , -4.332    , -4.685            // 3125
        , -4.508    , -4.862            // 3126
        , -4.508    , -4.685            // 3127
        , -4.862    , -4.332            // 3128
        , -4.862    , -4.508            // 3129
        , -4.685    , -4.332            // 3130
        , -4.685    , -4.508            // 3131
        , -4.862    , -4.862            // 3132
        , -4.862    , -4.685            // 3133
        , -4.685    , -4.862            // 3134
        , -4.685    , -4.685            // 3135
        , -5.569    , -2.917            // 3136
        , -5.569    , -3.094            // 3137
        , -5.392    , -2.917            // 3138
        , -5.392    , -3.094            // 3139
        , -5.569    , -3.448            // 3140
        , -5.569    , -3.271            // 3141
        , -5.392    , -3.448            // 3142
        , -5.392    , -3.271            // 3143
        , -5.039    , -2.917            // 3144
        , -5.039    , -3.094            // 3145
        , -5.216    , -2.917            // 3146
        , -5.216    , -3.094            // 3147
        , -5.039    , -3.448            // 3148
        , -5.039    , -3.271            // 3149
        , -5.216    , -3.448            // 3150
        , -5.216    , -3.271            // 3151
        , -5.569    , -4.155            // 3152
        , -5.569    , -3.978            // 3153
        , -5.392    , -4.155            // 3154
        , -5.392    , -3.978            // 3155
        , -5.569    , -3.624            // 3156
        , -5.569    , -3.801            // 3157
        , -5.392    , -3.624            // 3158
        , -5.392    , -3.801            // 3159
        , -5.039    , -4.155            // 3160
        , -5.039    , -3.978            // 3161
        , -5.216    , -4.155            // 3162
        , -5.216    , -3.978            // 3163
        , -5.039    , -3.624            // 3164
        , -5.039    , -3.801            // 3165
        , -5.216    , -3.624            // 3166
        , -5.216    , -3.801            // 3167
        , -4.332    , -2.917            // 3168
        , -4.332    , -3.094            // 3169
        , -4.508    , -2.917            // 3170
        , -4.508    , -3.094            // 3171
        , -4.332    , -3.448            // 3172
        , -4.332    , -3.271            // 3173
        , -4.508    , -3.448            // 3174
        , -4.508    , -3.271            // 3175
        , -4.862    , -2.917            // 3176
        , -4.862    , -3.094            // 3177
        , -4.685    , -2.917            // 3178
        , -4.685    , -3.094            // 3179
        , -4.862    , -3.448            // 3180
        , -4.862    , -3.271            // 3181
        , -4.685    , -3.448            // 3182
        , -4.685    , -3.271            // 3183
        , -4.332    , -4.155            // 3184
        , -4.332    , -3.978            // 3185
        , -4.508    , -4.155            // 3186
        , -4.508    , -3.978            // 3187
        , -4.332    , -3.624            // 3188
        , -4.332    , -3.801            // 3189
        , -4.508    , -3.624            // 3190
        , -4.508    , -3.801            // 3191
        , -4.862    , -4.155            // 3192
        , -4.862    , -3.978            // 3193
        , -4.685    , -4.155            // 3194
        , -4.685    , -3.978            // 3195
        , -4.862    , -3.624            // 3196
        , -4.862    , -3.801            // 3197
        , -4.685    , -3.624            // 3198
        , -4.685    , -3.801            // 3199
        , -2.917    , -5.569            // 3200
        , -2.917    , -5.392            // 3201
        , -3.094    , -5.569            // 3202
        , -3.094    , -5.392            // 3203
        , -2.917    , -5.039            // 3204
        , -2.917    , -5.216            // 3205
        , -3.094    , -5.039            // 3206
        , -3.094    , -5.216            // 3207
        , -3.448    , -5.569            // 3208
        , -3.448    , -5.392            // 3209
        , -3.271    , -5.569            // 3210
        , -3.271    , -5.392            // 3211
        , -3.448    , -5.039            // 3212
        , -3.448    , -5.216            // 3213
        , -3.271    , -5.039            // 3214
        , -3.271    , -5.216            // 3215
        , -2.917    , -4.332            // 3216
        , -2.917    , -4.508            // 3217
        , -3.094    , -4.332            // 3218
        , -3.094    , -4.508            // 3219
        , -2.917    , -4.862            // 3220
        , -2.917    , -4.685            // 3221
        , -3.094    , -4.862            // 3222
        , -3.094    , -4.685            // 3223
        , -3.448    , -4.332            // 3224
        , -3.448    , -4.508            // 3225
        , -3.271    , -4.332            // 3226
        , -3.271    , -4.508            // 3227
        , -3.448    , -4.862            // 3228
        , -3.448    , -4.685            // 3229
        , -3.271    , -4.862            // 3230
        , -3.271    , -4.685            // 3231
        , -4.155    , -5.569            // 3232
        , -4.155    , -5.392            // 3233
        , -3.978    , -5.569            // 3234
        , -3.978    , -5.392            // 3235
        , -4.155    , -5.039            // 3236
        , -4.155    , -5.216            // 3237
        , -3.978    , -5.039            // 3238
        , -3.978    , -5.216            // 3239
        , -3.624    , -5.569            // 3240
        , -3.624    , -5.392            // 3241
        , -3.801    , -5.569            // 3242
        , -3.801    , -5.392            // 3243
        , -3.624    , -5.039            // 3244
        , -3.624    , -5.216            // 3245
        , -3.801    , -5.039            // 3246
        , -3.801    , -5.216            // 3247
        , -4.155    , -4.332            // 3248
        , -4.155    , -4.508            // 3249
        , -3.978    , -4.332            // 3250
        , -3.978    , -4.508            // 3251
        , -4.155    , -4.862            // 3252
        , -4.155    , -4.685            // 3253
        , -3.978    , -4.862            // 3254
        , -3.978    , -4.685            // 3255
        , -3.624    , -4.332            // 3256
        , -3.624    , -4.508            // 3257
        , -3.801    , -4.332            // 3258
        , -3.801    , -4.508            // 3259
        , -3.624    , -4.862            // 3260
        , -3.624    , -4.685            // 3261
        , -3.801    , -4.862            // 3262
        , -3.801    , -4.685            // 3263
        , -2.917    , -2.917            // 3264
        , -2.917    , -3.094            // 3265
        , -3.094    , -2.917            // 3266
        , -3.094    , -3.094            // 3267
        , -2.917    , -3.448            // 3268
        , -2.917    , -3.271            // 3269
        , -3.094    , -3.448            // 3270
        , -3.094    , -3.271            // 3271
        , -3.448    , -2.917            // 3272
        , -3.448    , -3.094            // 3273
        , -3.271    , -2.917            // 3274
        , -3.271    , -3.094            // 3275
        , -3.448    , -3.448            // 3276
        , -3.448    , -3.271            // 3277
        , -3.271    , -3.448            // 3278
        , -3.271    , -3.271            // 3279
        , -2.917    , -4.155            // 3280
        , -2.917    , -3.978            // 3281
        , -3.094    , -4.155            // 3282
        , -3.094    , -3.978            // 3283
        , -2.917    , -3.624            // 3284
        , -2.917    , -3.801            // 3285
        , -3.094    , -3.624            // 3286
        , -3.094    , -3.801            // 3287
        , -3.448    , -4.155            // 3288
        , -3.448    , -3.978            // 3289
        , -3.271    , -4.155            // 3290
        , -3.271    , -3.978            // 3291
        , -3.448    , -3.624            // 3292
        , -3.448    , -3.801            // 3293
        , -3.271    , -3.624            // 3294
        , -3.271    , -3.801            // 3295
        , -4.155    , -2.917            // 3296
        , -4.155    , -3.094            // 3297
        , -3.978    , -2.917            // 3298
        , -3.978    , -3.094            // 3299
        , -4.155    , -3.448            // 3300
        , -4.155    , -3.271            // 3301
        , -3.978    , -3.448            // 3302
        , -3.978    , -3.271            // 3303
        , -3.624    , -2.917            // 3304
        , -3.624    , -3.094            // 3305
        , -3.801    , -2.917            // 3306
        , -3.801    , -3.094            // 3307
        , -3.624    , -3.448            // 3308
        , -3.624    , -3.271            // 3309
        , -3.801    , -3.448            // 3310
        , -3.801    , -3.271            // 3311
        , -4.155    , -4.155            // 3312
        , -4.155    , -3.978            // 3313
        , -3.978    , -4.155            // 3314
        , -3.978    , -3.978            // 3315
        , -4.155    , -3.624            // 3316
        , -4.155    , -3.801            // 3317
        , -3.978    , -3.624            // 3318
        , -3.978    , -3.801            // 3319
        , -3.624    , -4.155            // 3320
        , -3.624    , -3.978            // 3321
        , -3.801    , -4.155            // 3322
        , -3.801    , -3.978            // 3323
        , -3.624    , -3.624            // 3324
        , -3.624    , -3.801            // 3325
        , -3.801    , -3.624            // 3326
        , -3.801    , -3.801            // 3327
        , -5.569    , -0.088            // 3328
        , -5.569    , -0.265            // 3329
        , -5.392    , -0.088            // 3330
        , -5.392    , -0.265            // 3331
        , -5.569    , -0.619            // 3332
        , -5.569    , -0.442            // 3333
        , -5.392    , -0.619            // 3334
        , -5.392    , -0.442            // 3335
        , -5.039    , -0.088            // 3336
        , -5.039    , -0.265            // 3337
        , -5.216    , -0.088            // 3338
        , -5.216    , -0.265            // 3339
        , -5.039    , -0.619            // 3340
        , -5.039    , -0.442            // 3341
        , -5.216    , -0.619            // 3342
        , -5.216    , -0.442            // 3343
        , -5.569    , -1.326            // 3344
        , -5.569    , -1.149            // 3345
        , -5.392    , -1.326            // 3346
        , -5.392    , -1.149            // 3347
        , -5.569    , -0.796            // 3348
        , -5.569    , -0.972            // 3349
        , -5.392    , -0.796            // 3350
        , -5.392    , -0.972            // 3351
        , -5.039    , -1.326            // 3352
        , -5.039    , -1.149            // 3353
        , -5.216    , -1.326            // 3354
        , -5.216    , -1.149            // 3355
        , -5.039    , -0.796            // 3356
        , -5.039    , -0.972            // 3357
        , -5.216    , -0.796            // 3358
        , -5.216    , -0.972            // 3359
        , -4.332    , -0.088            // 3360
        , -4.332    , -0.265            // 3361
        , -4.508    , -0.088            // 3362
        , -4.508    , -0.265            // 3363
        , -4.332    , -0.619            // 3364
        , -4.332    , -0.442            // 3365
        , -4.508    , -0.619            // 3366
        , -4.508    , -0.442            // 3367
        , -4.862    , -0.088            // 3368
        , -4.862    , -0.265            // 3369
        , -4.685    , -0.088            // 3370
        , -4.685    , -0.265            // 3371
        , -4.862    , -0.619            // 3372
        , -4.862    , -0.442            // 3373
        , -4.685    , -0.619            // 3374
        , -4.685    , -0.442            // 3375
        , -4.332    , -1.326            // 3376
        , -4.332    , -1.149            // 3377
        , -4.508    , -1.326            // 3378
        , -4.508    , -1.149            // 3379
        , -4.332    , -0.796            // 3380
        , -4.332    , -0.972            // 3381
        , -4.508    , -0.796            // 3382
        , -4.508    , -0.972            // 3383
        , -4.862    , -1.326            // 3384
        , -4.862    , -1.149            // 3385
        , -4.685    , -1.326            // 3386
        , -4.685    , -1.149            // 3387
        , -4.862    , -0.796            // 3388
        , -4.862    , -0.972            // 3389
        , -4.685    , -0.796            // 3390
        , -4.685    , -0.972            // 3391
        , -5.569    ,  -2.74            // 3392
        , -5.569    , -2.564            // 3393
        , -5.392    ,  -2.74            // 3394
        , -5.392    , -2.564            // 3395
        , -5.569    ,  -2.21            // 3396
        , -5.569    , -2.387            // 3397
        , -5.392    ,  -2.21            // 3398
        , -5.392    , -2.387            // 3399
        , -5.039    ,  -2.74            // 3400
        , -5.039    , -2.564            // 3401
        , -5.216    ,  -2.74            // 3402
        , -5.216    , -2.564            // 3403
        , -5.039    ,  -2.21            // 3404
        , -5.039    , -2.387            // 3405
        , -5.216    ,  -2.21            // 3406
        , -5.216    , -2.387            // 3407
        , -5.569    , -1.503            // 3408
        , -5.569    ,  -1.68            // 3409
        , -5.392    , -1.503            // 3410
        , -5.392    ,  -1.68            // 3411
        , -5.569    , -2.033            // 3412
        , -5.569    , -1.856            // 3413
        , -5.392    , -2.033            // 3414
        , -5.392    , -1.856            // 3415
        , -5.039    , -1.503            // 3416
        , -5.039    ,  -1.68            // 3417
        , -5.216    , -1.503            // 3418
        , -5.216    ,  -1.68            // 3419
        , -5.039    , -2.033            // 3420
        , -5.039    , -1.856            // 3421
        , -5.216    , -2.033            // 3422
        , -5.216    , -1.856            // 3423
        , -4.332    ,  -2.74            // 3424
        , -4.332    , -2.564            // 3425
        , -4.508    ,  -2.74            // 3426
        , -4.508    , -2.564            // 3427
        , -4.332    ,  -2.21            // 3428
        , -4.332    , -2.387            // 3429
        , -4.508    ,  -2.21            // 3430
        , -4.508    , -2.387            // 3431
        , -4.862    ,  -2.74            // 3432
        , -4.862    , -2.564            // 3433
        , -4.685    ,  -2.74            // 3434
        , -4.685    , -2.564            // 3435
        , -4.862    ,  -2.21            // 3436
        , -4.862    , -2.387            // 3437
        , -4.685    ,  -2.21            // 3438
        , -4.685    , -2.387            // 3439
        , -4.332    , -1.503            // 3440
        , -4.332    ,  -1.68            // 3441
        , -4.508    , -1.503            // 3442
        , -4.508    ,  -1.68            // 3443
        , -4.332    , -2.033            // 3444
        , -4.332    , -1.856            // 3445
        , -4.508    , -2.033            // 3446
        , -4.508    , -1.856            // 3447
        , -4.862    , -1.503            // 3448
        , -4.862    ,  -1.68            // 3449
        , -4.685    , -1.503            // 3450
        , -4.685    ,  -1.68            // 3451
        , -4.862    , -2.033            // 3452
        , -4.862    , -1.856            // 3453
        , -4.685    , -2.033            // 3454
        , -4.685    , -1.856            // 3455
        , -2.917    , -0.088            // 3456
        , -2.917    , -0.265            // 3457
        , -3.094    , -0.088            // 3458
        , -3.094    , -0.265            // 3459
        , -2.917    , -0.619            // 3460
        , -2.917    , -0.442            // 3461
        , -3.094    , -0.619            // 3462
        , -3.094    , -0.442            // 3463
        , -3.448    , -0.088            // 3464
        , -3.448    , -0.265            // 3465
        , -3.271    , -0.088            // 3466
        , -3.271    , -0.265            // 3467
        , -3.448    , -0.619            // 3468
        , -3.448    , -0.442            // 3469
        , -3.271    , -0.619            // 3470
        , -3.271    , -0.442            // 3471
        , -2.917    , -1.326            // 3472
        , -2.917    , -1.149            // 3473
        , -3.094    , -1.326            // 3474
        , -3.094    , -1.149            // 3475
        , -2.917    , -0.796            // 3476
        , -2.917    , -0.972            // 3477
        , -3.094    , -0.796            // 3478
        , -3.094    , -0.972            // 3479
        , -3.448    , -1.326            // 3480
        , -3.448    , -1.149            // 3481
        , -3.271    , -1.326            // 3482
        , -3.271    , -1.149            // 3483
        , -3.448    , -0.796            // 3484
        , -3.448    , -0.972            // 3485
        , -3.271    , -0.796            // 3486
        , -3.271    , -0.972            // 3487
        , -4.155    , -0.088            // 3488
        , -4.155    , -0.265            // 3489
        , -3.978    , -0.088            // 3490
        , -3.978    , -0.265            // 3491
        , -4.155    , -0.619            // 3492
        , -4.155    , -0.442            // 3493
        , -3.978    , -0.619            // 3494
        , -3.978    , -0.442            // 3495
        , -3.624    , -0.088            // 3496
        , -3.624    , -0.265            // 3497
        , -3.801    , -0.088            // 3498
        , -3.801    , -0.265            // 3499
        , -3.624    , -0.619            // 3500
        , -3.624    , -0.442            // 3501
        , -3.801    , -0.619            // 3502
        , -3.801    , -0.442            // 3503
        , -4.155    , -1.326            // 3504
        , -4.155    , -1.149            // 3505
        , -3.978    , -1.326            // 3506
        , -3.978    , -1.149            // 3507
        , -4.155    , -0.796            // 3508
        , -4.155    , -0.972            // 3509
        , -3.978    , -0.796            // 3510
        , -3.978    , -0.972            // 3511
        , -3.624    , -1.326            // 3512
        , -3.624    , -1.149            // 3513
        , -3.801    , -1.326            // 3514
        , -3.801    , -1.149            // 3515
        , -3.624    , -0.796            // 3516
        , -3.624    , -0.972            // 3517
        , -3.801    , -0.796            // 3518
        , -3.801    , -0.972            // 3519
        , -2.917    ,  -2.74            // 3520
        , -2.917    , -2.564            // 3521
        , -3.094    ,  -2.74            // 3522
        , -3.094    , -2.564            // 3523
        , -2.917    ,  -2.21            // 3524
        , -2.917    , -2.387            // 3525
        , -3.094    ,  -2.21            // 3526
        , -3.094    , -2.387            // 3527
        , -3.448    ,  -2.74            // 3528
        , -3.448    , -2.564            // 3529
        , -3.271    ,  -2.74            // 3530
        , -3.271    , -2.564            // 3531
        , -3.448    ,  -2.21            // 3532
        , -3.448    , -2.387            // 3533
        , -3.271    ,  -2.21            // 3534
        , -3.271    , -2.387            // 3535
        , -2.917    , -1.503            // 3536
        , -2.917    ,  -1.68            // 3537
        , -3.094    , -1.503            // 3538
        , -3.094    ,  -1.68            // 3539
        , -2.917    , -2.033            // 3540
        , -2.917    , -1.856            // 3541
        , -3.094    , -2.033            // 3542
        , -3.094    , -1.856            // 3543
        , -3.448    , -1.503            // 3544
        , -3.448    ,  -1.68            // 3545
        , -3.271    , -1.503            // 3546
        , -3.271    ,  -1.68            // 3547
        , -3.448    , -2.033            // 3548
        , -3.448    , -1.856            // 3549
        , -3.271    , -2.033            // 3550
        , -3.271    , -1.856            // 3551
        , -4.155    ,  -2.74            // 3552
        , -4.155    , -2.564            // 3553
        , -3.978    ,  -2.74            // 3554
        , -3.978    , -2.564            // 3555
        , -4.155    ,  -2.21            // 3556
        , -4.155    , -2.387            // 3557
        , -3.978    ,  -2.21            // 3558
        , -3.978    , -2.387            // 3559
        , -3.624    ,  -2.74            // 3560
        , -3.624    , -2.564            // 3561
        , -3.801    ,  -2.74            // 3562
        , -3.801    , -2.564            // 3563
        , -3.624    ,  -2.21            // 3564
        , -3.624    , -2.387            // 3565
        , -3.801    ,  -2.21            // 3566
        , -3.801    , -2.387            // 3567
        , -4.155    , -1.503            // 3568
        , -4.155    ,  -1.68            // 3569
        , -3.978    , -1.503            // 3570
        , -3.978    ,  -1.68            // 3571
        , -4.155    , -2.033            // 3572
        , -4.155    , -1.856            // 3573
        , -3.978    , -2.033            // 3574
        , -3.978    , -1.856            // 3575
        , -3.624    , -1.503            // 3576
        , -3.624    ,  -1.68            // 3577
        , -3.801    , -1.503            // 3578
        , -3.801    ,  -1.68            // 3579
        , -3.624    , -2.033            // 3580
        , -3.624    , -1.856            // 3581
        , -3.801    , -2.033            // 3582
        , -3.801    , -1.856            // 3583
        , -0.088    , -5.569            // 3584
        , -0.088    , -5.392            // 3585
        , -0.265    , -5.569            // 3586
        , -0.265    , -5.392            // 3587
        , -0.088    , -5.039            // 3588
        , -0.088    , -5.216            // 3589
        , -0.265    , -5.039            // 3590
        , -0.265    , -5.216            // 3591
        , -0.619    , -5.569            // 3592
        , -0.619    , -5.392            // 3593
        , -0.442    , -5.569            // 3594
        , -0.442    , -5.392            // 3595
        , -0.619    , -5.039            // 3596
        , -0.619    , -5.216            // 3597
        , -0.442    , -5.039            // 3598
        , -0.442    , -5.216            // 3599
        , -0.088    , -4.332            // 3600
        , -0.088    , -4.508            // 3601
        , -0.265    , -4.332            // 3602
        , -0.265    , -4.508            // 3603
        , -0.088    , -4.862            // 3604
        , -0.088    , -4.685            // 3605
        , -0.265    , -4.862            // 3606
        , -0.265    , -4.685            // 3607
        , -0.619    , -4.332            // 3608
        , -0.619    , -4.508            // 3609
        , -0.442    , -4.332            // 3610
        , -0.442    , -4.508            // 3611
        , -0.619    , -4.862            // 3612
        , -0.619    , -4.685            // 3613
        , -0.442    , -4.862            // 3614
        , -0.442    , -4.685            // 3615
        , -1.326    , -5.569            // 3616
        , -1.326    , -5.392            // 3617
        , -1.149    , -5.569            // 3618
        , -1.149    , -5.392            // 3619
        , -1.326    , -5.039            // 3620
        , -1.326    , -5.216            // 3621
        , -1.149    , -5.039            // 3622
        , -1.149    , -5.216            // 3623
        , -0.796    , -5.569            // 3624
        , -0.796    , -5.392            // 3625
        , -0.972    , -5.569            // 3626
        , -0.972    , -5.392            // 3627
        , -0.796    , -5.039            // 3628
        , -0.796    , -5.216            // 3629
        , -0.972    , -5.039            // 3630
        , -0.972    , -5.216            // 3631
        , -1.326    , -4.332            // 3632
        , -1.326    , -4.508            // 3633
        , -1.149    , -4.332            // 3634
        , -1.149    , -4.508            // 3635
        , -1.326    , -4.862            // 3636
        , -1.326    , -4.685            // 3637
        , -1.149    , -4.862            // 3638
        , -1.149    , -4.685            // 3639
        , -0.796    , -4.332            // 3640
        , -0.796    , -4.508            // 3641
        , -0.972    , -4.332            // 3642
        , -0.972    , -4.508            // 3643
        , -0.796    , -4.862            // 3644
        , -0.796    , -4.685            // 3645
        , -0.972    , -4.862            // 3646
        , -0.972    , -4.685            // 3647
        , -0.088    , -2.917            // 3648
        , -0.088    , -3.094            // 3649
        , -0.265    , -2.917            // 3650
        , -0.265    , -3.094            // 3651
        , -0.088    , -3.448            // 3652
        , -0.088    , -3.271            // 3653
        , -0.265    , -3.448            // 3654
        , -0.265    , -3.271            // 3655
        , -0.619    , -2.917            // 3656
        , -0.619    , -3.094            // 3657
        , -0.442    , -2.917            // 3658
        , -0.442    , -3.094            // 3659
        , -0.619    , -3.448            // 3660
        , -0.619    , -3.271            // 3661
        , -0.442    , -3.448            // 3662
        , -0.442    , -3.271            // 3663
        , -0.088    , -4.155            // 3664
        , -0.088    , -3.978            // 3665
        , -0.265    , -4.155            // 3666
        , -0.265    , -3.978            // 3667
        , -0.088    , -3.624            // 3668
        , -0.088    , -3.801            // 3669
        , -0.265    , -3.624            // 3670
        , -0.265    , -3.801            // 3671
        , -0.619    , -4.155            // 3672
        , -0.619    , -3.978            // 3673
        , -0.442    , -4.155            // 3674
        , -0.442    , -3.978            // 3675
        , -0.619    , -3.624            // 3676
        , -0.619    , -3.801            // 3677
        , -0.442    , -3.624            // 3678
        , -0.442    , -3.801            // 3679
        , -1.326    , -2.917            // 3680
        , -1.326    , -3.094            // 3681
        , -1.149    , -2.917            // 3682
        , -1.149    , -3.094            // 3683
        , -1.326    , -3.448            // 3684
        , -1.326    , -3.271            // 3685
        , -1.149    , -3.448            // 3686
        , -1.149    , -3.271            // 3687
        , -0.796    , -2.917            // 3688
        , -0.796    , -3.094            // 3689
        , -0.972    , -2.917            // 3690
        , -0.972    , -3.094            // 3691
        , -0.796    , -3.448            // 3692
        , -0.796    , -3.271            // 3693
        , -0.972    , -3.448            // 3694
        , -0.972    , -3.271            // 3695
        , -1.326    , -4.155            // 3696
        , -1.326    , -3.978            // 3697
        , -1.149    , -4.155            // 3698
        , -1.149    , -3.978            // 3699
        , -1.326    , -3.624            // 3700
        , -1.326    , -3.801            // 3701
        , -1.149    , -3.624            // 3702
        , -1.149    , -3.801            // 3703
        , -0.796    , -4.155            // 3704
        , -0.796    , -3.978            // 3705
        , -0.972    , -4.155            // 3706
        , -0.972    , -3.978            // 3707
        , -0.796    , -3.624            // 3708
        , -0.796    , -3.801            // 3709
        , -0.972    , -3.624            // 3710
        , -0.972    , -3.801            // 3711
        ,  -2.74    , -5.569            // 3712
        ,  -2.74    , -5.392            // 3713
        , -2.564    , -5.569            // 3714
        , -2.564    , -5.392            // 3715
        ,  -2.74    , -5.039            // 3716
        ,  -2.74    , -5.216            // 3717
        , -2.564    , -5.039            // 3718
        , -2.564    , -5.216            // 3719
        ,  -2.21    , -5.569            // 3720
        ,  -2.21    , -5.392            // 3721
        , -2.387    , -5.569            // 3722
        , -2.387    , -5.392            // 3723
        ,  -2.21    , -5.039            // 3724
        ,  -2.21    , -5.216            // 3725
        , -2.387    , -5.039            // 3726
        , -2.387    , -5.216            // 3727
        ,  -2.74    , -4.332            // 3728
        ,  -2.74    , -4.508            // 3729
        , -2.564    , -4.332            // 3730
        , -2.564    , -4.508            // 3731
        ,  -2.74    , -4.862            // 3732
        ,  -2.74    , -4.685            // 3733
        , -2.564    , -4.862            // 3734
        , -2.564    , -4.685            // 3735
        ,  -2.21    , -4.332            // 3736
        ,  -2.21    , -4.508            // 3737
        , -2.387    , -4.332            // 3738
        , -2.387    , -4.508            // 3739
        ,  -2.21    , -4.862            // 3740
        ,  -2.21    , -4.685            // 3741
        , -2.387    , -4.862            // 3742
        , -2.387    , -4.685            // 3743
        , -1.503    , -5.569            // 3744
        , -1.503    , -5.392            // 3745
        ,  -1.68    , -5.569            // 3746
        ,  -1.68    , -5.392            // 3747
        , -1.503    , -5.039            // 3748
        , -1.503    , -5.216            // 3749
        ,  -1.68    , -5.039            // 3750
        ,  -1.68    , -5.216            // 3751
        , -2.033    , -5.569            // 3752
        , -2.033    , -5.392            // 3753
        , -1.856    , -5.569            // 3754
        , -1.856    , -5.392            // 3755
        , -2.033    , -5.039            // 3756
        , -2.033    , -5.216            // 3757
        , -1.856    , -5.039            // 3758
        , -1.856    , -5.216            // 3759
        , -1.503    , -4.332            // 3760
        , -1.503    , -4.508            // 3761
        ,  -1.68    , -4.332            // 3762
        ,  -1.68    , -4.508            // 3763
        , -1.503    , -4.862            // 3764
        , -1.503    , -4.685            // 3765
        ,  -1.68    , -4.862            // 3766
        ,  -1.68    , -4.685            // 3767
        , -2.033    , -4.332            // 3768
        , -2.033    , -4.508            // 3769
        , -1.856    , -4.332            // 3770
        , -1.856    , -4.508            // 3771
        , -2.033    , -4.862            // 3772
        , -2.033    , -4.685            // 3773
        , -1.856    , -4.862            // 3774
        , -1.856    , -4.685            // 3775
        ,  -2.74    , -2.917            // 3776
        ,  -2.74    , -3.094            // 3777
        , -2.564    , -2.917            // 3778
        , -2.564    , -3.094            // 3779
        ,  -2.74    , -3.448            // 3780
        ,  -2.74    , -3.271            // 3781
        , -2.564    , -3.448            // 3782
        , -2.564    , -3.271            // 3783
        ,  -2.21    , -2.917            // 3784
        ,  -2.21    , -3.094            // 3785
        , -2.387    , -2.917            // 3786
        , -2.387    , -3.094            // 3787
        ,  -2.21    , -3.448            // 3788
        ,  -2.21    , -3.271            // 3789
        , -2.387    , -3.448            // 3790
        , -2.387    , -3.271            // 3791
        ,  -2.74    , -4.155            // 3792
        ,  -2.74    , -3.978            // 3793
        , -2.564    , -4.155            // 3794
        , -2.564    , -3.978            // 3795
        ,  -2.74    , -3.624            // 3796
        ,  -2.74    , -3.801            // 3797
        , -2.564    , -3.624            // 3798
        , -2.564    , -3.801            // 3799
        ,  -2.21    , -4.155            // 3800
        ,  -2.21    , -3.978            // 3801
        , -2.387    , -4.155            // 3802
        , -2.387    , -3.978            // 3803
        ,  -2.21    , -3.624            // 3804
        ,  -2.21    , -3.801            // 3805
        , -2.387    , -3.624            // 3806
        , -2.387    , -3.801            // 3807
        , -1.503    , -2.917            // 3808
        , -1.503    , -3.094            // 3809
        ,  -1.68    , -2.917            // 3810
        ,  -1.68    , -3.094            // 3811
        , -1.503    , -3.448            // 3812
        , -1.503    , -3.271            // 3813
        ,  -1.68    , -3.448            // 3814
        ,  -1.68    , -3.271            // 3815
        , -2.033    , -2.917            // 3816
        , -2.033    , -3.094            // 3817
        , -1.856    , -2.917            // 3818
        , -1.856    , -3.094            // 3819
        , -2.033    , -3.448            // 3820
        , -2.033    , -3.271            // 3821
        , -1.856    , -3.448            // 3822
        , -1.856    , -3.271            // 3823
        , -1.503    , -4.155            // 3824
        , -1.503    , -3.978            // 3825
        ,  -1.68    , -4.155            // 3826
        ,  -1.68    , -3.978            // 3827
        , -1.503    , -3.624            // 3828
        , -1.503    , -3.801            // 3829
        ,  -1.68    , -3.624            // 3830
        ,  -1.68    , -3.801            // 3831
        , -2.033    , -4.155            // 3832
        , -2.033    , -3.978            // 3833
        , -1.856    , -4.155            // 3834
        , -1.856    , -3.978            // 3835
        , -2.033    , -3.624            // 3836
        , -2.033    , -3.801            // 3837
        , -1.856    , -3.624            // 3838
        , -1.856    , -3.801            // 3839
        , -0.088    , -0.088            // 3840
        , -0.088    , -0.265            // 3841
        , -0.265    , -0.088            // 3842
        , -0.265    , -0.265            // 3843
        , -0.088    , -0.619            // 3844
        , -0.088    , -0.442            // 3845
        , -0.265    , -0.619            // 3846
        , -0.265    , -0.442            // 3847
        , -0.619    , -0.088            // 3848
        , -0.619    , -0.265            // 3849
        , -0.442    , -0.088            // 3850
        , -0.442    , -0.265            // 3851
        , -0.619    , -0.619            // 3852
        , -0.619    , -0.442            // 3853
        , -0.442    , -0.619            // 3854
        , -0.442    , -0.442            // 3855
        , -0.088    , -1.326            // 3856
        , -0.088    , -1.149            // 3857
        , -0.265    , -1.326            // 3858
        , -0.265    , -1.149            // 3859
        , -0.088    , -0.796            // 3860
        , -0.088    , -0.972            // 3861
        , -0.265    , -0.796            // 3862
        , -0.265    , -0.972            // 3863
        , -0.619    , -1.326            // 3864
        , -0.619    , -1.149            // 3865
        , -0.442    , -1.326            // 3866
        , -0.442    , -1.149            // 3867
        , -0.619    , -0.796            // 3868
        , -0.619    , -0.972            // 3869
        , -0.442    , -0.796            // 3870
        , -0.442    , -0.972            // 3871
        , -1.326    , -0.088            // 3872
        , -1.326    , -0.265            // 3873
        , -1.149    , -0.088            // 3874
        , -1.149    , -0.265            // 3875
        , -1.326    , -0.619            // 3876
        , -1.326    , -0.442            // 3877
        , -1.149    , -0.619            // 3878
        , -1.149    , -0.442            // 3879
        , -0.796    , -0.088            // 3880
        , -0.796    , -0.265            // 3881
        , -0.972    , -0.088            // 3882
        , -0.972    , -0.265            // 3883
        , -0.796    , -0.619            // 3884
        , -0.796    , -0.442            // 3885
        , -0.972    , -0.619            // 3886
        , -0.972    , -0.442            // 3887
        , -1.326    , -1.326            // 3888
        , -1.326    , -1.149            // 3889
        , -1.149    , -1.326            // 3890
        , -1.149    , -1.149            // 3891
        , -1.326    , -0.796            // 3892
        , -1.326    , -0.972            // 3893
        , -1.149    , -0.796            // 3894
        , -1.149    , -0.972            // 3895
        , -0.796    , -1.326            // 3896
        , -0.796    , -1.149            // 3897
        , -0.972    , -1.326            // 3898
        , -0.972    , -1.149            // 3899
        , -0.796    , -0.796            // 3900
        , -0.796    , -0.972            // 3901
        , -0.972    , -0.796            // 3902
        , -0.972    , -0.972            // 3903
        , -0.088    ,  -2.74            // 3904
        , -0.088    , -2.564            // 3905
        , -0.265    ,  -2.74            // 3906
        , -0.265    , -2.564            // 3907
        , -0.088    ,  -2.21            // 3908
        , -0.088    , -2.387            // 3909
        , -0.265    ,  -2.21            // 3910
        , -0.265    , -2.387            // 3911
        , -0.619    ,  -2.74            // 3912
        , -0.619    , -2.564            // 3913
        , -0.442    ,  -2.74            // 3914
        , -0.442    , -2.564            // 3915
        , -0.619    ,  -2.21            // 3916
        , -0.619    , -2.387            // 3917
        , -0.442    ,  -2.21            // 3918
        , -0.442    , -2.387            // 3919
        , -0.088    , -1.503            // 3920
        , -0.088    ,  -1.68            // 3921
        , -0.265    , -1.503            // 3922
        , -0.265    ,  -1.68            // 3923
        , -0.088    , -2.033            // 3924
        , -0.088    , -1.856            // 3925
        , -0.265    , -2.033            // 3926
        , -0.265    , -1.856            // 3927
        , -0.619    , -1.503            // 3928
        , -0.619    ,  -1.68            // 3929
        , -0.442    , -1.503            // 3930
        , -0.442    ,  -1.68            // 3931
        , -0.619    , -2.033            // 3932
        , -0.619    , -1.856            // 3933
        , -0.442    , -2.033            // 3934
        , -0.442    , -1.856            // 3935
        , -1.326    ,  -2.74            // 3936
        , -1.326    , -2.564            // 3937
        , -1.149    ,  -2.74            // 3938
        , -1.149    , -2.564            // 3939
        , -1.326    ,  -2.21            // 3940
        , -1.326    , -2.387            // 3941
        , -1.149    ,  -2.21            // 3942
        , -1.149    , -2.387            // 3943
        , -0.796    ,  -2.74            // 3944
        , -0.796    , -2.564            // 3945
        , -0.972    ,  -2.74            // 3946
        , -0.972    , -2.564            // 3947
        , -0.796    ,  -2.21            // 3948
        , -0.796    , -2.387            // 3949
        , -0.972    ,  -2.21            // 3950
        , -0.972    , -2.387            // 3951
        , -1.326    , -1.503            // 3952
        , -1.326    ,  -1.68            // 3953
        , -1.149    , -1.503            // 3954
        , -1.149    ,  -1.68            // 3955
        , -1.326    , -2.033            // 3956
        , -1.326    , -1.856            // 3957
        , -1.149    , -2.033            // 3958
        , -1.149    , -1.856            // 3959
        , -0.796    , -1.503            // 3960
        , -0.796    ,  -1.68            // 3961
        , -0.972    , -1.503            // 3962
        , -0.972    ,  -1.68            // 3963
        , -0.796    , -2.033            // 3964
        , -0.796    , -1.856            // 3965
        , -0.972    , -2.033            // 3966
        , -0.972    , -1.856            // 3967
        ,  -2.74    , -0.088            // 3968
        ,  -2.74    , -0.265            // 3969
        , -2.564    , -0.088            // 3970
        , -2.564    , -0.265            // 3971
        ,  -2.74    , -0.619            // 3972
        ,  -2.74    , -0.442            // 3973
        , -2.564    , -0.619            // 3974
        , -2.564    , -0.442            // 3975
        ,  -2.21    , -0.088            // 3976
        ,  -2.21    , -0.265            // 3977
        , -2.387    , -0.088            // 3978
        , -2.387    , -0.265            // 3979
        ,  -2.21    , -0.619            // 3980
        ,  -2.21    , -0.442            // 3981
        , -2.387    , -0.619            // 3982
        , -2.387    , -0.442            // 3983
        ,  -2.74    , -1.326            // 3984
        ,  -2.74    , -1.149            // 3985
        , -2.564    , -1.326            // 3986
        , -2.564    , -1.149            // 3987
        ,  -2.74    , -0.796            // 3988
        ,  -2.74    , -0.972            // 3989
        , -2.564    , -0.796            // 3990
        , -2.564    , -0.972            // 3991
        ,  -2.21    , -1.326            // 3992
        ,  -2.21    , -1.149            // 3993
        , -2.387    , -1.326            // 3994
        , -2.387    , -1.149            // 3995
        ,  -2.21    , -0.796            // 3996
        ,  -2.21    , -0.972            // 3997
        , -2.387    , -0.796            // 3998
        , -2.387    , -0.972            // 3999
        , -1.503    , -0.088            // 4000
        , -1.503    , -0.265            // 4001
        ,  -1.68    , -0.088            // 4002
        ,  -1.68    , -0.265            // 4003
        , -1.503    , -0.619            // 4004
        , -1.503    , -0.442            // 4005
        ,  -1.68    , -0.619            // 4006
        ,  -1.68    , -0.442            // 4007
        , -2.033    , -0.088            // 4008
        , -2.033    , -0.265            // 4009
        , -1.856    , -0.088            // 4010
        , -1.856    , -0.265            // 4011
        , -2.033    , -0.619            // 4012
        , -2.033    , -0.442            // 4013
        , -1.856    , -0.619            // 4014
        , -1.856    , -0.442            // 4015
        , -1.503    , -1.326            // 4016
        , -1.503    , -1.149            // 4017
        ,  -1.68    , -1.326            // 4018
        ,  -1.68    , -1.149            // 4019
        , -1.503    , -0.796            // 4020
        , -1.503    , -0.972            // 4021
        ,  -1.68    , -0.796            // 4022
        ,  -1.68    , -0.972            // 4023
        , -2.033    , -1.326            // 4024
        , -2.033    , -1.149            // 4025
        , -1.856    , -1.326            // 4026
        , -1.856    , -1.149            // 4027
        , -2.033    , -0.796            // 4028
        , -2.033    , -0.972            // 4029
        , -1.856    , -0.796            // 4030
        , -1.856    , -0.972            // 4031
        ,  -2.74    ,  -2.74            // 4032
        ,  -2.74    , -2.564            // 4033
        , -2.564    ,  -2.74            // 4034
        , -2.564    , -2.564            // 4035
        ,  -2.74    ,  -2.21            // 4036
        ,  -2.74    , -2.387            // 4037
        , -2.564    ,  -2.21            // 4038
        , -2.564    , -2.387            // 4039
        ,  -2.21    ,  -2.74            // 4040
        ,  -2.21    , -2.564            // 4041
        , -2.387    ,  -2.74            // 4042
        , -2.387    , -2.564            // 4043
        ,  -2.21    ,  -2.21            // 4044
        ,  -2.21    , -2.387            // 4045
        , -2.387    ,  -2.21            // 4046
        , -2.387    , -2.387            // 4047
        ,  -2.74    , -1.503            // 4048
        ,  -2.74    ,  -1.68            // 4049
        , -2.564    , -1.503            // 4050
        , -2.564    ,  -1.68            // 4051
        ,  -2.74    , -2.033            // 4052
        ,  -2.74    , -1.856            // 4053
        , -2.564    , -2.033            // 4054
        , -2.564    , -1.856            // 4055
        ,  -2.21    , -1.503            // 4056
        ,  -2.21    ,  -1.68            // 4057
        , -2.387    , -1.503            // 4058
        , -2.387    ,  -1.68            // 4059
        ,  -2.21    , -2.033            // 4060
        ,  -2.21    , -1.856            // 4061
        , -2.387    , -2.033            // 4062
        , -2.387    , -1.856            // 4063
        , -1.503    ,  -2.74            // 4064
        , -1.503    , -2.564            // 4065
        ,  -1.68    ,  -2.74            // 4066
        ,  -1.68    , -2.564            // 4067
        , -1.503    ,  -2.21            // 4068
        , -1.503    , -2.387            // 4069
        ,  -1.68    ,  -2.21            // 4070
        ,  -1.68    , -2.387            // 4071
        , -2.033    ,  -2.74            // 4072
        , -2.033    , -2.564            // 4073
        , -1.856    ,  -2.74            // 4074
        , -1.856    , -2.564            // 4075
        , -2.033    ,  -2.21            // 4076
        , -2.033    , -2.387            // 4077
        , -1.856    ,  -2.21            // 4078
        , -1.856    , -2.387            // 4079
        , -1.503    , -1.503            // 4080
        , -1.503    ,  -1.68            // 4081
        ,  -1.68    , -1.503            // 4082
        ,  -1.68    ,  -1.68            // 4083
        , -1.503    , -2.033            // 4084
        , -1.503    , -1.856            // 4085
        ,  -1.68    , -2.033            // 4086
        ,  -1.68    , -1.856            // 4087
        , -2.033    , -1.503            // 4088
        , -2.033    ,  -1.68            // 4089
        , -1.856    , -1.503            // 4090
        , -1.856    ,  -1.68            // 4091
        , -2.033    , -2.033            // 4092
        , -2.033    , -1.856            // 4093
        , -1.856    , -2.033            // 4094
        , -1.856    , -1.856            // 4095
    };