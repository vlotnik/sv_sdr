    DVBS2X_256APSK_20_30 : super.plane = {
           1.635    ,  0.159            // 0
        ,  1.578    ,  0.474            // 1
        ,  0.943    ,   0.11            // 2
        ,  0.907    ,  0.283            // 3
        ,  0.324    ,  0.085            // 4
        ,  0.323    ,  0.087            // 5
        ,   0.75    ,  0.114            // 6
        ,  0.733    ,  0.209            // 7
        ,  0.166    ,  1.675            // 8
        ,  0.491    ,  1.608            // 9
        ,  0.109    ,  0.953            // 10
        ,  0.246    ,  0.927            // 11
        ,  0.087    ,  0.139            // 12
        ,  0.087    ,  0.139            // 13
        ,  0.109    ,  0.766            // 14
        ,   0.17    ,  0.754            // 15
        , -1.635    ,  0.159            // 16
        , -1.578    ,  0.474            // 17
        , -0.943    ,   0.11            // 18
        , -0.907    ,  0.283            // 19
        , -0.324    ,  0.085            // 20
        , -0.323    ,  0.087            // 21
        ,  -0.75    ,  0.114            // 22
        , -0.733    ,  0.209            // 23
        , -0.166    ,  1.675            // 24
        , -0.491    ,  1.608            // 25
        , -0.109    ,  0.953            // 26
        , -0.246    ,  0.927            // 27
        , -0.087    ,  0.139            // 28
        , -0.087    ,  0.139            // 29
        , -0.109    ,  0.766            // 30
        ,  -0.17    ,  0.754            // 31
        ,  1.323    ,  0.132            // 32
        ,  1.274    ,  0.392            // 33
        ,  1.085    ,  0.114            // 34
        ,  1.044    ,   0.33            // 35
        ,  0.458    ,  0.112            // 36
        ,  0.455    ,  0.125            // 37
        ,  0.647    ,  0.114            // 38
        ,  0.634    ,   0.17            // 39
        ,  0.132    ,  1.363            // 40
        ,  0.393    ,   1.31            // 41
        ,  0.112    ,  1.133            // 42
        ,  0.316    ,  1.091            // 43
        ,  0.093    ,  0.397            // 44
        ,  0.094    ,  0.397            // 45
        ,  0.105    ,  0.598            // 46
        ,  0.123    ,  0.595            // 47
        , -1.323    ,  0.132            // 48
        , -1.274    ,  0.392            // 49
        , -1.085    ,  0.114            // 50
        , -1.044    ,   0.33            // 51
        , -0.458    ,  0.112            // 52
        , -0.455    ,  0.125            // 53
        , -0.647    ,  0.114            // 54
        , -0.634    ,   0.17            // 55
        , -0.132    ,  1.363            // 56
        , -0.393    ,   1.31            // 57
        , -0.112    ,  1.133            // 58
        , -0.316    ,  1.091            // 59
        , -0.093    ,  0.397            // 60
        , -0.094    ,  0.397            // 61
        , -0.105    ,  0.598            // 62
        , -0.123    ,  0.595            // 63
        ,  1.635    , -0.159            // 64
        ,  1.578    , -0.474            // 65
        ,  0.943    ,  -0.11            // 66
        ,  0.907    , -0.283            // 67
        ,  0.324    , -0.085            // 68
        ,  0.323    , -0.087            // 69
        ,   0.75    , -0.114            // 70
        ,  0.733    , -0.209            // 71
        ,  0.166    , -1.675            // 72
        ,  0.491    , -1.608            // 73
        ,  0.109    , -0.953            // 74
        ,  0.246    , -0.927            // 75
        ,  0.087    , -0.139            // 76
        ,  0.087    , -0.139            // 77
        ,  0.109    , -0.766            // 78
        ,   0.17    , -0.754            // 79
        , -1.635    , -0.159            // 80
        , -1.578    , -0.474            // 81
        , -0.943    ,  -0.11            // 82
        , -0.907    , -0.283            // 83
        , -0.324    , -0.085            // 84
        , -0.323    , -0.087            // 85
        ,  -0.75    , -0.114            // 86
        , -0.733    , -0.209            // 87
        , -0.166    , -1.675            // 88
        , -0.491    , -1.608            // 89
        , -0.109    , -0.953            // 90
        , -0.246    , -0.927            // 91
        , -0.087    , -0.139            // 92
        , -0.087    , -0.139            // 93
        , -0.109    , -0.766            // 94
        ,  -0.17    , -0.754            // 95
        ,  1.323    , -0.132            // 96
        ,  1.274    , -0.392            // 97
        ,  1.085    , -0.114            // 98
        ,  1.044    ,  -0.33            // 99
        ,  0.458    , -0.112            // 100
        ,  0.455    , -0.125            // 101
        ,  0.647    , -0.114            // 102
        ,  0.634    ,  -0.17            // 103
        ,  0.132    , -1.363            // 104
        ,  0.393    ,  -1.31            // 105
        ,  0.112    , -1.133            // 106
        ,  0.316    , -1.091            // 107
        ,  0.093    , -0.397            // 108
        ,  0.094    , -0.397            // 109
        ,  0.105    , -0.598            // 110
        ,  0.123    , -0.595            // 111
        , -1.323    , -0.132            // 112
        , -1.274    , -0.392            // 113
        , -1.085    , -0.114            // 114
        , -1.044    ,  -0.33            // 115
        , -0.458    , -0.112            // 116
        , -0.455    , -0.125            // 117
        , -0.647    , -0.114            // 118
        , -0.634    ,  -0.17            // 119
        , -0.132    , -1.363            // 120
        , -0.393    ,  -1.31            // 121
        , -0.112    , -1.133            // 122
        , -0.316    , -1.091            // 123
        , -0.093    , -0.397            // 124
        , -0.094    , -0.397            // 125
        , -0.105    , -0.598            // 126
        , -0.123    , -0.595            // 127
        ,   1.29    ,   1.05            // 128
        ,  1.463    ,  0.774            // 129
        ,  0.727    ,  0.616            // 130
        ,  0.818    ,  0.484            // 131
        ,  0.284    ,   0.13            // 132
        ,  0.285    ,  0.131            // 133
        ,   0.59    ,  0.486            // 134
        ,  0.636    ,  0.419            // 135
        ,  1.065    ,  1.288            // 136
        ,  0.795    ,  1.477            // 137
        ,  0.571    ,  0.766            // 138
        ,  0.449    ,  0.846            // 139
        ,  0.105    ,  0.149            // 140
        ,  0.105    ,   0.15            // 141
        ,  0.429    ,  0.636            // 142
        ,  0.374    ,  0.674            // 143
        ,  -1.29    ,   1.05            // 144
        , -1.463    ,  0.774            // 145
        , -0.727    ,  0.616            // 146
        , -0.818    ,  0.484            // 147
        , -0.284    ,   0.13            // 148
        , -0.285    ,  0.131            // 149
        ,  -0.59    ,  0.486            // 150
        , -0.636    ,  0.419            // 151
        , -1.065    ,  1.288            // 152
        , -0.795    ,  1.477            // 153
        , -0.571    ,  0.766            // 154
        , -0.449    ,  0.846            // 155
        , -0.105    ,  0.149            // 156
        , -0.105    ,   0.15            // 157
        , -0.429    ,  0.636            // 158
        , -0.374    ,  0.674            // 159
        ,  1.038    ,  0.862            // 160
        ,  1.179    ,  0.638            // 161
        ,   0.85    ,  0.722            // 162
        ,  0.964    ,  0.541            // 163
        ,  0.373    ,  0.256            // 164
        ,   0.38    ,  0.252            // 165
        ,  0.497    ,  0.395            // 166
        ,  0.523    ,  0.364            // 167
        ,  0.856    ,  1.054            // 168
        ,  0.636    ,  1.206            // 169
        ,  0.696    ,  0.885            // 170
        ,  0.523    ,  1.004            // 171
        ,  0.194    ,  0.362            // 172
        ,  0.191    ,  0.363            // 173
        ,  0.322    ,  0.524            // 174
        ,  0.302    ,  0.535            // 175
        , -1.038    ,  0.862            // 176
        , -1.179    ,  0.638            // 177
        ,  -0.85    ,  0.722            // 178
        , -0.964    ,  0.541            // 179
        , -0.373    ,  0.256            // 180
        ,  -0.38    ,  0.252            // 181
        , -0.497    ,  0.395            // 182
        , -0.523    ,  0.364            // 183
        , -0.856    ,  1.054            // 184
        , -0.636    ,  1.206            // 185
        , -0.696    ,  0.885            // 186
        , -0.523    ,  1.004            // 187
        , -0.194    ,  0.362            // 188
        , -0.191    ,  0.363            // 189
        , -0.322    ,  0.524            // 190
        , -0.302    ,  0.535            // 191
        ,   1.29    ,  -1.05            // 192
        ,  1.463    , -0.774            // 193
        ,  0.727    , -0.616            // 194
        ,  0.818    , -0.484            // 195
        ,  0.284    ,  -0.13            // 196
        ,  0.285    , -0.131            // 197
        ,   0.59    , -0.486            // 198
        ,  0.636    , -0.419            // 199
        ,  1.065    , -1.288            // 200
        ,  0.795    , -1.477            // 201
        ,  0.571    , -0.766            // 202
        ,  0.449    , -0.846            // 203
        ,  0.105    , -0.149            // 204
        ,  0.105    ,  -0.15            // 205
        ,  0.429    , -0.636            // 206
        ,  0.374    , -0.674            // 207
        ,  -1.29    ,  -1.05            // 208
        , -1.463    , -0.774            // 209
        , -0.727    , -0.616            // 210
        , -0.818    , -0.484            // 211
        , -0.284    ,  -0.13            // 212
        , -0.285    , -0.131            // 213
        ,  -0.59    , -0.486            // 214
        , -0.636    , -0.419            // 215
        , -1.065    , -1.288            // 216
        , -0.795    , -1.477            // 217
        , -0.571    , -0.766            // 218
        , -0.449    , -0.846            // 219
        , -0.105    , -0.149            // 220
        , -0.105    ,  -0.15            // 221
        , -0.429    , -0.636            // 222
        , -0.374    , -0.674            // 223
        ,  1.038    , -0.862            // 224
        ,  1.179    , -0.638            // 225
        ,   0.85    , -0.722            // 226
        ,  0.964    , -0.541            // 227
        ,  0.373    , -0.256            // 228
        ,   0.38    , -0.252            // 229
        ,  0.497    , -0.395            // 230
        ,  0.523    , -0.364            // 231
        ,  0.856    , -1.054            // 232
        ,  0.636    , -1.206            // 233
        ,  0.696    , -0.885            // 234
        ,  0.523    , -1.004            // 235
        ,  0.194    , -0.362            // 236
        ,  0.191    , -0.363            // 237
        ,  0.322    , -0.524            // 238
        ,  0.302    , -0.535            // 239
        , -1.038    , -0.862            // 240
        , -1.179    , -0.638            // 241
        ,  -0.85    , -0.722            // 242
        , -0.964    , -0.541            // 243
        , -0.373    , -0.256            // 244
        ,  -0.38    , -0.252            // 245
        , -0.497    , -0.395            // 246
        , -0.523    , -0.364            // 247
        , -0.856    , -1.054            // 248
        , -0.636    , -1.206            // 249
        , -0.696    , -0.885            // 250
        , -0.523    , -1.004            // 251
        , -0.194    , -0.362            // 252
        , -0.191    , -0.363            // 253
        , -0.322    , -0.524            // 254
        , -0.302    , -0.535            // 255
    };