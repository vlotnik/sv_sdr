    DVBS2_APSK16_2_3 : super.plane = {
           0.803    ,  0.803            // 0
        ,  0.803    , -0.803            // 1
        , -0.803    ,  0.803            // 2
        , -0.803    , -0.803            // 3
        ,  1.097    ,  0.294            // 4
        ,  1.097    , -0.294            // 5
        , -1.097    ,  0.294            // 6
        , -1.097    , -0.294            // 7
        ,  0.294    ,  1.097            // 8
        ,  0.294    , -1.097            // 9
        , -0.294    ,  1.097            // 10
        , -0.294    , -1.097            // 11
        ,  0.255    ,  0.255            // 12
        ,  0.255    , -0.255            // 13
        , -0.255    ,  0.255            // 14
        , -0.255    , -0.255            // 15
    };