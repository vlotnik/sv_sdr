    QAM32 : super.plane = {
            1.33    ,  0.798            // 0
        ,  0.798    ,  0.798            // 1
        ,  0.798    ,   1.33            // 2
        ,  0.798    ,  0.266            // 3
        ,   1.33    ,  0.266            // 4
        ,  0.266    ,  0.798            // 5
        ,  0.266    ,   1.33            // 6
        ,  0.266    ,  0.266            // 7
        ,  0.798    ,  -1.33            // 8
        ,  0.798    , -0.798            // 9
        ,   1.33    , -0.798            // 10
        ,  0.266    , -0.798            // 11
        ,  0.266    ,  -1.33            // 12
        ,  0.798    , -0.266            // 13
        ,   1.33    , -0.266            // 14
        ,  0.266    , -0.266            // 15
        , -0.798    ,   1.33            // 16
        , -0.798    ,  0.798            // 17
        ,  -1.33    ,  0.798            // 18
        , -0.266    ,  0.798            // 19
        , -0.266    ,   1.33            // 20
        , -0.798    ,  0.266            // 21
        ,  -1.33    ,  0.266            // 22
        , -0.266    ,  0.266            // 23
        ,  -1.33    , -0.798            // 24
        , -0.798    , -0.798            // 25
        , -0.798    ,  -1.33            // 26
        , -0.798    , -0.266            // 27
        ,  -1.33    , -0.266            // 28
        , -0.266    , -0.798            // 29
        , -0.266    ,  -1.33            // 30
        , -0.266    , -0.266            // 31
    };