    DVBS2X_APSK8_L_5_9 : super.plane = {
          -0.196    ,      0            // 0
        , -0.468    , -0.934            // 1
        , -0.468    ,  0.934            // 2
        , -1.335    ,      0            // 3
        ,  0.196    ,      0            // 4
        ,  0.468    , -0.934            // 5
        ,  0.468    ,  0.934            // 6
        ,  1.335    ,      0            // 7
    };