    DVBS2X_8_8APSK_18_30 : super.plane = {
           0.472    ,  0.261            // 0
        ,  0.261    ,  0.472            // 1
        , -0.472    ,  0.261            // 2
        , -0.261    ,  0.472            // 3
        ,  0.472    , -0.261            // 4
        ,  0.261    , -0.472            // 5
        , -0.472    , -0.261            // 6
        , -0.261    , -0.472            // 7
        ,  1.209    ,  0.498            // 8
        ,  0.498    ,  1.209            // 9
        , -1.209    ,  0.498            // 10
        , -0.498    ,  1.209            // 11
        ,  1.209    , -0.498            // 12
        ,  0.498    , -1.209            // 13
        , -1.209    , -0.498            // 14
        , -0.498    , -1.209            // 15
    };