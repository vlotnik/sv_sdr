    DVBS2_QPSK : super.plane = {
           0.707    ,  0.707            // 0
        ,  0.707    , -0.707            // 1
        , -0.707    ,  0.707            // 2
        , -0.707    , -0.707            // 3
    };