    PSK8 : super.plane = {
           1.000    ,  0.000            // 0
        ,  0.707    ,  0.707            // 1
        ,  0.000    ,  1.000            // 2
        , -0.707    ,  0.707            // 3
        , -1.000    ,  0.000            // 4
        , -0.707    , -0.707            // 5
        ,  0.000    , -1.000            // 6
        ,  0.707    , -0.707            // 7
    };