    DVBS2X_8_16_20_20APSK_4_5 : super.plane = {
           0.115    ,  -0.58            // 0
        ,  0.989    , -0.989            // 1
        ,  0.329    , -0.492            // 2
        ,  0.685    , -0.685            // 3
        ,  0.219    , -1.382            // 4
        ,  0.635    , -1.246            // 5
        ,  0.151    , -0.956            // 6
        ,   0.44    , -0.863            // 7
        , -0.115    ,  -0.58            // 8
        , -0.989    , -0.989            // 9
        , -0.329    , -0.492            // 10
        , -0.685    , -0.685            // 11
        , -0.219    , -1.382            // 12
        , -0.635    , -1.246            // 13
        , -0.151    , -0.956            // 14
        ,  -0.44    , -0.863            // 15
        ,  0.103    , -0.249            // 16
        ,  1.246    , -0.635            // 17
        ,  0.492    , -0.329            // 18
        ,  0.863    ,  -0.44            // 19
        ,  0.249    , -0.103            // 20
        ,  1.382    , -0.219            // 21
        ,   0.58    , -0.115            // 22
        ,  0.956    , -0.151            // 23
        , -0.103    , -0.249            // 24
        , -1.246    , -0.635            // 25
        , -0.492    , -0.329            // 26
        , -0.863    ,  -0.44            // 27
        , -0.249    , -0.103            // 28
        , -1.382    , -0.219            // 29
        ,  -0.58    , -0.115            // 30
        , -0.956    , -0.151            // 31
        ,  0.115    ,   0.58            // 32
        ,  0.989    ,  0.989            // 33
        ,  0.329    ,  0.492            // 34
        ,  0.685    ,  0.685            // 35
        ,  0.219    ,  1.382            // 36
        ,  0.635    ,  1.246            // 37
        ,  0.151    ,  0.956            // 38
        ,   0.44    ,  0.863            // 39
        , -0.115    ,   0.58            // 40
        , -0.989    ,  0.989            // 41
        , -0.329    ,  0.492            // 42
        , -0.685    ,  0.685            // 43
        , -0.219    ,  1.382            // 44
        , -0.635    ,  1.246            // 45
        , -0.151    ,  0.956            // 46
        ,  -0.44    ,  0.863            // 47
        ,  0.103    ,  0.249            // 48
        ,  1.246    ,  0.635            // 49
        ,  0.492    ,  0.329            // 50
        ,  0.863    ,   0.44            // 51
        ,  0.249    ,  0.103            // 52
        ,  1.382    ,  0.219            // 53
        ,   0.58    ,  0.115            // 54
        ,  0.956    ,  0.151            // 55
        , -0.103    ,  0.249            // 56
        , -1.246    ,  0.635            // 57
        , -0.492    ,  0.329            // 58
        , -0.863    ,   0.44            // 59
        , -0.249    ,  0.103            // 60
        , -1.382    ,  0.219            // 61
        ,  -0.58    ,  0.115            // 62
        , -0.956    ,  0.151            // 63
    };