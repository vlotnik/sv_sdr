    DVBS2_APSK16_8_9 : super.plane = {
           0.797    ,  0.797            // 0
        ,  0.797    , -0.797            // 1
        , -0.797    ,  0.797            // 2
        , -0.797    , -0.797            // 3
        ,  1.089    ,  0.292            // 4
        ,  1.089    , -0.292            // 5
        , -1.089    ,  0.292            // 6
        , -1.089    , -0.292            // 7
        ,  0.292    ,  1.089            // 8
        ,  0.292    , -1.089            // 9
        , -0.292    ,  1.089            // 10
        , -0.292    , -1.089            // 11
        ,  0.307    ,  0.307            // 12
        ,  0.307    , -0.307            // 13
        , -0.307    ,  0.307            // 14
        , -0.307    , -0.307            // 15
    };