    DVBS2X_256APSK_128_180 : super.plane = {
           0.284    ,  0.028            // 0
        ,  0.273    ,  0.083            // 1
        ,   0.22    ,  0.181            // 2
        ,  0.251    ,  0.134            // 3
        ,  0.028    ,  0.284            // 4
        ,  0.083    ,  0.273            // 5
        ,  0.181    ,   0.22            // 6
        ,  0.134    ,  0.251            // 7
        , -0.284    ,  0.028            // 8
        , -0.273    ,  0.083            // 9
        ,  -0.22    ,  0.181            // 10
        , -0.251    ,  0.134            // 11
        , -0.028    ,  0.284            // 12
        , -0.083    ,  0.273            // 13
        , -0.181    ,   0.22            // 14
        , -0.134    ,  0.251            // 15
        ,  0.284    , -0.028            // 16
        ,  0.273    , -0.083            // 17
        ,   0.22    , -0.181            // 18
        ,  0.251    , -0.134            // 19
        ,  0.028    , -0.284            // 20
        ,  0.083    , -0.273            // 21
        ,  0.181    ,  -0.22            // 22
        ,  0.134    , -0.251            // 23
        , -0.284    , -0.028            // 24
        , -0.273    , -0.083            // 25
        ,  -0.22    , -0.181            // 26
        , -0.251    , -0.134            // 27
        , -0.028    , -0.284            // 28
        , -0.083    , -0.273            // 29
        , -0.181    ,  -0.22            // 30
        , -0.134    , -0.251            // 31
        ,  0.509    ,   0.05            // 32
        ,  0.489    ,  0.148            // 33
        ,  0.395    ,  0.324            // 34
        ,  0.451    ,  0.241            // 35
        ,   0.05    ,  0.509            // 36
        ,  0.148    ,  0.489            // 37
        ,  0.324    ,  0.395            // 38
        ,  0.241    ,  0.451            // 39
        , -0.509    ,   0.05            // 40
        , -0.489    ,  0.148            // 41
        , -0.395    ,  0.324            // 42
        , -0.451    ,  0.241            // 43
        ,  -0.05    ,  0.509            // 44
        , -0.148    ,  0.489            // 45
        , -0.324    ,  0.395            // 46
        , -0.241    ,  0.451            // 47
        ,  0.509    ,  -0.05            // 48
        ,  0.489    , -0.148            // 49
        ,  0.395    , -0.324            // 50
        ,  0.451    , -0.241            // 51
        ,   0.05    , -0.509            // 52
        ,  0.148    , -0.489            // 53
        ,  0.324    , -0.395            // 54
        ,  0.241    , -0.451            // 55
        , -0.509    ,  -0.05            // 56
        , -0.489    , -0.148            // 57
        , -0.395    , -0.324            // 58
        , -0.451    , -0.241            // 59
        ,  -0.05    , -0.509            // 60
        , -0.148    , -0.489            // 61
        , -0.324    , -0.395            // 62
        , -0.241    , -0.451            // 63
        ,  0.847    ,  0.083            // 64
        ,  0.815    ,  0.247            // 65
        ,  0.658    ,   0.54            // 66
        ,  0.751    ,  0.401            // 67
        ,  0.083    ,  0.847            // 68
        ,  0.247    ,  0.815            // 69
        ,   0.54    ,  0.658            // 70
        ,  0.401    ,  0.751            // 71
        , -0.847    ,  0.083            // 72
        , -0.815    ,  0.247            // 73
        , -0.658    ,   0.54            // 74
        , -0.751    ,  0.401            // 75
        , -0.083    ,  0.847            // 76
        , -0.247    ,  0.815            // 77
        ,  -0.54    ,  0.658            // 78
        , -0.401    ,  0.751            // 79
        ,  0.847    , -0.083            // 80
        ,  0.815    , -0.247            // 81
        ,  0.658    ,  -0.54            // 82
        ,  0.751    , -0.401            // 83
        ,  0.083    , -0.847            // 84
        ,  0.247    , -0.815            // 85
        ,   0.54    , -0.658            // 86
        ,  0.401    , -0.751            // 87
        , -0.847    , -0.083            // 88
        , -0.815    , -0.247            // 89
        , -0.658    ,  -0.54            // 90
        , -0.751    , -0.401            // 91
        , -0.083    , -0.847            // 92
        , -0.247    , -0.815            // 93
        ,  -0.54    , -0.658            // 94
        , -0.401    , -0.751            // 95
        ,  0.683    ,  0.067            // 96
        ,  0.657    ,  0.199            // 97
        ,  0.531    ,  0.436            // 98
        ,  0.606    ,  0.324            // 99
        ,  0.067    ,  0.683            // 100
        ,  0.199    ,  0.657            // 101
        ,  0.436    ,  0.531            // 102
        ,  0.324    ,  0.606            // 103
        , -0.683    ,  0.067            // 104
        , -0.657    ,  0.199            // 105
        , -0.531    ,  0.436            // 106
        , -0.606    ,  0.324            // 107
        , -0.067    ,  0.683            // 108
        , -0.199    ,  0.657            // 109
        , -0.436    ,  0.531            // 110
        , -0.324    ,  0.606            // 111
        ,  0.683    , -0.067            // 112
        ,  0.657    , -0.199            // 113
        ,  0.531    , -0.436            // 114
        ,  0.606    , -0.324            // 115
        ,  0.067    , -0.683            // 116
        ,  0.199    , -0.657            // 117
        ,  0.436    , -0.531            // 118
        ,  0.324    , -0.606            // 119
        , -0.683    , -0.067            // 120
        , -0.657    , -0.199            // 121
        , -0.531    , -0.436            // 122
        , -0.606    , -0.324            // 123
        , -0.067    , -0.683            // 124
        , -0.199    , -0.657            // 125
        , -0.436    , -0.531            // 126
        , -0.324    , -0.606            // 127
        ,  1.532    ,  0.151            // 128
        ,  1.473    ,  0.447            // 129
        ,   1.19    ,  0.977            // 130
        ,  1.358    ,  0.726            // 131
        ,  0.151    ,  1.532            // 132
        ,  0.447    ,  1.473            // 133
        ,  0.977    ,   1.19            // 134
        ,  0.726    ,  1.358            // 135
        , -1.532    ,  0.151            // 136
        , -1.473    ,  0.447            // 137
        ,  -1.19    ,  0.977            // 138
        , -1.358    ,  0.726            // 139
        , -0.151    ,  1.532            // 140
        , -0.447    ,  1.473            // 141
        , -0.977    ,   1.19            // 142
        , -0.726    ,  1.358            // 143
        ,  1.532    , -0.151            // 144
        ,  1.473    , -0.447            // 145
        ,   1.19    , -0.977            // 146
        ,  1.358    , -0.726            // 147
        ,  0.151    , -1.532            // 148
        ,  0.447    , -1.473            // 149
        ,  0.977    ,  -1.19            // 150
        ,  0.726    , -1.358            // 151
        , -1.532    , -0.151            // 152
        , -1.473    , -0.447            // 153
        ,  -1.19    , -0.977            // 154
        , -1.358    , -0.726            // 155
        , -0.151    , -1.532            // 156
        , -0.447    , -1.473            // 157
        , -0.977    ,  -1.19            // 158
        , -0.726    , -1.358            // 159
        ,  1.305    ,  0.129            // 160
        ,  1.255    ,  0.381            // 161
        ,  1.014    ,  0.832            // 162
        ,  1.157    ,  0.618            // 163
        ,  0.129    ,  1.305            // 164
        ,  0.381    ,  1.255            // 165
        ,  0.832    ,  1.014            // 166
        ,  0.618    ,  1.157            // 167
        , -1.305    ,  0.129            // 168
        , -1.255    ,  0.381            // 169
        , -1.014    ,  0.832            // 170
        , -1.157    ,  0.618            // 171
        , -0.129    ,  1.305            // 172
        , -0.381    ,  1.255            // 173
        , -0.832    ,  1.014            // 174
        , -0.618    ,  1.157            // 175
        ,  1.305    , -0.129            // 176
        ,  1.255    , -0.381            // 177
        ,  1.014    , -0.832            // 178
        ,  1.157    , -0.618            // 179
        ,  0.129    , -1.305            // 180
        ,  0.381    , -1.255            // 181
        ,  0.832    , -1.014            // 182
        ,  0.618    , -1.157            // 183
        , -1.305    , -0.129            // 184
        , -1.255    , -0.381            // 185
        , -1.014    , -0.832            // 186
        , -1.157    , -0.618            // 187
        , -0.129    , -1.305            // 188
        , -0.381    , -1.255            // 189
        , -0.832    , -1.014            // 190
        , -0.618    , -1.157            // 191
        ,  1.015    ,    0.1            // 192
        ,  0.976    ,  0.296            // 193
        ,  0.789    ,  0.647            // 194
        ,    0.9    ,  0.481            // 195
        ,    0.1    ,  1.015            // 196
        ,  0.296    ,  0.976            // 197
        ,  0.647    ,  0.789            // 198
        ,  0.481    ,    0.9            // 199
        , -1.015    ,    0.1            // 200
        , -0.976    ,  0.296            // 201
        , -0.789    ,  0.647            // 202
        ,   -0.9    ,  0.481            // 203
        ,   -0.1    ,  1.015            // 204
        , -0.296    ,  0.976            // 205
        , -0.647    ,  0.789            // 206
        , -0.481    ,    0.9            // 207
        ,  1.015    ,   -0.1            // 208
        ,  0.976    , -0.296            // 209
        ,  0.789    , -0.647            // 210
        ,    0.9    , -0.481            // 211
        ,    0.1    , -1.015            // 212
        ,  0.296    , -0.976            // 213
        ,  0.647    , -0.789            // 214
        ,  0.481    ,   -0.9            // 215
        , -1.015    ,   -0.1            // 216
        , -0.976    , -0.296            // 217
        , -0.789    , -0.647            // 218
        ,   -0.9    , -0.481            // 219
        ,   -0.1    , -1.015            // 220
        , -0.296    , -0.976            // 221
        , -0.647    , -0.789            // 222
        , -0.481    ,   -0.9            // 223
        ,  1.148    ,  0.113            // 224
        ,  1.104    ,  0.335            // 225
        ,  0.891    ,  0.732            // 226
        ,  1.017    ,  0.544            // 227
        ,  0.113    ,  1.148            // 228
        ,  0.335    ,  1.104            // 229
        ,  0.732    ,  0.891            // 230
        ,  0.544    ,  1.017            // 231
        , -1.148    ,  0.113            // 232
        , -1.104    ,  0.335            // 233
        , -0.891    ,  0.732            // 234
        , -1.017    ,  0.544            // 235
        , -0.113    ,  1.148            // 236
        , -0.335    ,  1.104            // 237
        , -0.732    ,  0.891            // 238
        , -0.544    ,  1.017            // 239
        ,  1.148    , -0.113            // 240
        ,  1.104    , -0.335            // 241
        ,  0.891    , -0.732            // 242
        ,  1.017    , -0.544            // 243
        ,  0.113    , -1.148            // 244
        ,  0.335    , -1.104            // 245
        ,  0.732    , -0.891            // 246
        ,  0.544    , -1.017            // 247
        , -1.148    , -0.113            // 248
        , -1.104    , -0.335            // 249
        , -0.891    , -0.732            // 250
        , -1.017    , -0.544            // 251
        , -0.113    , -1.148            // 252
        , -0.335    , -1.104            // 253
        , -0.732    , -0.891            // 254
        , -0.544    , -1.017            // 255
    };