    DVBS2_PSK8 : super.plane = {
           0.707    ,  0.707            // 0
        ,  1.000    ,  0.000            // 1
        , -1.000    ,  0.000            // 2
        , -0.707    , -0.707            // 3
        ,  0.000    ,  1.000            // 4
        ,  0.707    , -0.707            // 5
        , -0.707    ,  0.707            // 6
        ,  0.000    , -1.000            // 7
    };