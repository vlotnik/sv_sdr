    DVBS2X_4_8_4_16APSK_132_180 : super.plane = {
           0.164    ,  0.164            // 0
        ,  0.254    ,  1.277            // 1
        ,  0.164    , -0.164            // 2
        ,  0.254    , -1.277            // 3
        , -0.164    ,  0.164            // 4
        , -0.254    ,  1.277            // 5
        , -0.164    , -0.164            // 6
        , -0.254    , -1.277            // 7
        ,  0.584    ,  0.156            // 8
        ,  1.277    ,  0.254            // 9
        ,  0.584    , -0.156            // 10
        ,  1.277    , -0.254            // 11
        , -0.584    ,  0.156            // 12
        , -1.277    ,  0.254            // 13
        , -0.584    , -0.156            // 14
        , -1.277    , -0.254            // 15
        ,  0.156    ,  0.584            // 16
        ,  0.723    ,  1.083            // 17
        ,  0.156    , -0.584            // 18
        ,  0.723    , -1.083            // 19
        , -0.156    ,  0.584            // 20
        , -0.723    ,  1.083            // 21
        , -0.156    , -0.584            // 22
        , -0.723    , -1.083            // 23
        ,   0.47    ,   0.47            // 24
        ,  1.083    ,  0.723            // 25
        ,   0.47    ,  -0.47            // 26
        ,  1.083    , -0.723            // 27
        ,  -0.47    ,   0.47            // 28
        , -1.083    ,  0.723            // 29
        ,  -0.47    ,  -0.47            // 30
        , -1.083    , -0.723            // 31
    };