    DVBS2X_128APSK_140_180 : super.plane = {
           0.344    ,  0.072            // 0
        ,   1.24    ,  0.423            // 1
        ,  1.307    ,  0.091            // 2
        ,  1.283    ,  0.268            // 3
        ,  0.595    ,   0.09            // 4
        ,  0.719    ,   0.19            // 5
        ,  0.962    ,   0.08            // 6
        ,  0.908    ,  0.248            // 7
        ,  0.294    ,  0.192            // 8
        ,  1.176    ,  0.577            // 9
        ,  0.988    ,   0.86            // 10
        ,  1.097    ,  0.717            // 11
        ,  0.485    ,  0.357            // 12
        ,  0.643    ,  0.374            // 13
        ,  0.737    ,  0.623            // 14
        ,  0.817    ,  0.467            // 15
        ,  0.072    ,  0.343            // 16
        ,  0.423    ,   1.24            // 17
        ,  0.091    ,  1.307            // 18
        ,  0.268    ,  1.283            // 19
        ,   0.09    ,  0.595            // 20
        ,   0.19    ,  0.719            // 21
        ,   0.08    ,  0.962            // 22
        ,  0.247    ,  0.908            // 23
        ,  0.192    ,  0.294            // 24
        ,  0.577    ,  1.177            // 25
        ,   0.86    ,  0.989            // 26
        ,  0.718    ,  1.096            // 27
        ,  0.357    ,  0.485            // 28
        ,  0.375    ,  0.642            // 29
        ,  0.624    ,  0.737            // 30
        ,  0.467    ,  0.817            // 31
        , -0.344    ,  0.072            // 32
        ,  -1.24    ,  0.423            // 33
        , -1.307    ,  0.091            // 34
        , -1.283    ,  0.268            // 35
        , -0.595    ,   0.09            // 36
        , -0.719    ,   0.19            // 37
        , -0.962    ,   0.08            // 38
        , -0.908    ,  0.248            // 39
        , -0.294    ,  0.192            // 40
        , -1.176    ,  0.577            // 41
        , -0.988    ,   0.86            // 42
        , -1.097    ,  0.717            // 43
        , -0.485    ,  0.357            // 44
        , -0.643    ,  0.374            // 45
        , -0.737    ,  0.623            // 46
        , -0.817    ,  0.467            // 47
        , -0.072    ,  0.343            // 48
        , -0.423    ,   1.24            // 49
        , -0.091    ,  1.307            // 50
        , -0.268    ,  1.283            // 51
        ,  -0.09    ,  0.595            // 52
        ,  -0.19    ,  0.719            // 53
        ,  -0.08    ,  0.962            // 54
        , -0.247    ,  0.908            // 55
        , -0.192    ,  0.294            // 56
        , -0.577    ,  1.177            // 57
        ,  -0.86    ,  0.989            // 58
        , -0.718    ,  1.096            // 59
        , -0.357    ,  0.485            // 60
        , -0.375    ,  0.642            // 61
        , -0.624    ,  0.737            // 62
        , -0.467    ,  0.817            // 63
        ,  0.344    , -0.072            // 64
        ,   1.24    , -0.423            // 65
        ,  1.307    , -0.091            // 66
        ,  1.283    , -0.268            // 67
        ,  0.595    ,  -0.09            // 68
        ,  0.719    ,  -0.19            // 69
        ,  0.962    ,  -0.08            // 70
        ,  0.908    , -0.248            // 71
        ,  0.294    , -0.192            // 72
        ,  1.176    , -0.577            // 73
        ,  0.988    ,  -0.86            // 74
        ,  1.097    , -0.717            // 75
        ,  0.485    , -0.357            // 76
        ,  0.643    , -0.374            // 77
        ,  0.737    , -0.623            // 78
        ,  0.817    , -0.467            // 79
        ,  0.072    , -0.343            // 80
        ,  0.423    ,  -1.24            // 81
        ,  0.091    , -1.307            // 82
        ,  0.268    , -1.283            // 83
        ,   0.09    , -0.595            // 84
        ,   0.19    , -0.719            // 85
        ,   0.08    , -0.962            // 86
        ,  0.247    , -0.908            // 87
        ,  0.192    , -0.294            // 88
        ,  0.577    , -1.177            // 89
        ,   0.86    , -0.989            // 90
        ,  0.718    , -1.096            // 91
        ,  0.357    , -0.485            // 92
        ,  0.375    , -0.642            // 93
        ,  0.624    , -0.737            // 94
        ,  0.467    , -0.817            // 95
        , -0.344    , -0.072            // 96
        ,  -1.24    , -0.423            // 97
        , -1.307    , -0.091            // 98
        , -1.283    , -0.268            // 99
        , -0.595    ,  -0.09            // 100
        , -0.719    ,  -0.19            // 101
        , -0.962    ,  -0.08            // 102
        , -0.908    , -0.248            // 103
        , -0.294    , -0.192            // 104
        , -1.176    , -0.577            // 105
        , -0.988    ,  -0.86            // 106
        , -1.097    , -0.717            // 107
        , -0.485    , -0.357            // 108
        , -0.643    , -0.374            // 109
        , -0.737    , -0.623            // 110
        , -0.817    , -0.467            // 111
        , -0.072    , -0.343            // 112
        , -0.423    ,  -1.24            // 113
        , -0.091    , -1.307            // 114
        , -0.268    , -1.283            // 115
        ,  -0.09    , -0.595            // 116
        ,  -0.19    , -0.719            // 117
        ,  -0.08    , -0.962            // 118
        , -0.247    , -0.908            // 119
        , -0.192    , -0.294            // 120
        , -0.577    , -1.177            // 121
        ,  -0.86    , -0.989            // 122
        , -0.718    , -1.096            // 123
        , -0.357    , -0.485            // 124
        , -0.375    , -0.642            // 125
        , -0.624    , -0.737            // 126
        , -0.467    , -0.817            // 127
    };