    DVBS2X_4_12APSK_154_180 : super.plane = {
           0.804    ,  0.804            // 0
        ,  0.804    , -0.804            // 1
        , -0.804    ,  0.804            // 2
        , -0.804    , -0.804            // 3
        ,  1.098    ,  0.294            // 4
        ,  1.098    , -0.294            // 5
        , -1.098    ,  0.294            // 6
        , -1.098    , -0.294            // 7
        ,  0.294    ,  1.098            // 8
        ,  0.294    , -1.098            // 9
        , -0.294    ,  1.098            // 10
        , -0.294    , -1.098            // 11
        ,  0.251    ,  0.251            // 12
        ,  0.251    , -0.251            // 13
        , -0.251    ,  0.251            // 14
        , -0.251    , -0.251            // 15
    };