    DVBS2X_256APSK_22_30 : super.plane = {
           1.598    ,  0.153            // 0
        ,  1.319    ,  0.127            // 1
        , -1.598    ,  0.153            // 2
        , -1.319    ,  0.127            // 3
        ,  0.257    ,  0.073            // 4
        ,   0.45    ,  0.081            // 5
        , -0.257    ,  0.073            // 6
        ,  -0.45    ,  0.081            // 7
        ,  1.598    , -0.153            // 8
        ,  1.319    , -0.127            // 9
        , -1.598    , -0.153            // 10
        , -1.319    , -0.127            // 11
        ,  0.257    , -0.073            // 12
        ,   0.45    , -0.081            // 13
        , -0.257    , -0.073            // 14
        ,  -0.45    , -0.081            // 15
        ,  0.927    ,  0.094            // 16
        ,  1.102    ,  0.109            // 17
        , -0.927    ,  0.094            // 18
        , -1.102    ,  0.109            // 19
        ,  0.766    ,  0.087            // 20
        ,  0.612    ,  0.087            // 21
        , -0.766    ,  0.087            // 22
        , -0.612    ,  0.087            // 23
        ,  0.927    , -0.094            // 24
        ,  1.102    , -0.109            // 25
        , -0.927    , -0.094            // 26
        , -1.102    , -0.109            // 27
        ,  0.766    , -0.087            // 28
        ,  0.612    , -0.087            // 29
        , -0.766    , -0.087            // 30
        , -0.612    , -0.087            // 31
        ,   1.27    ,  1.014            // 32
        ,  1.053    ,  0.841            // 33
        ,  -1.27    ,  1.014            // 34
        , -1.053    ,  0.841            // 35
        ,  0.249    ,  0.198            // 36
        ,  0.352    ,  0.292            // 37
        , -0.249    ,  0.198            // 38
        , -0.352    ,  0.292            // 39
        ,   1.27    , -1.014            // 40
        ,  1.053    , -0.841            // 41
        ,  -1.27    , -1.014            // 42
        , -1.053    , -0.841            // 43
        ,  0.249    , -0.198            // 44
        ,  0.352    , -0.292            // 45
        , -0.249    , -0.198            // 46
        , -0.352    , -0.292            // 47
        ,  0.736    ,  0.604            // 48
        ,  0.881    ,  0.711            // 49
        , -0.736    ,  0.604            // 50
        , -0.881    ,  0.711            // 51
        ,  0.602    ,  0.502            // 52
        ,  0.475    ,    0.4            // 53
        , -0.602    ,  0.502            // 54
        , -0.475    ,    0.4            // 55
        ,  0.736    , -0.604            // 56
        ,  0.881    , -0.711            // 57
        , -0.736    , -0.604            // 58
        , -0.881    , -0.711            // 59
        ,  0.602    , -0.502            // 60
        ,  0.475    ,   -0.4            // 61
        , -0.602    , -0.502            // 62
        , -0.475    ,   -0.4            // 63
        ,  1.544    ,  0.455            // 64
        ,  1.275    ,  0.378            // 65
        , -1.544    ,  0.455            // 66
        , -1.275    ,  0.378            // 67
        ,  0.259    ,  0.075            // 68
        ,  0.444    ,  0.107            // 69
        , -0.259    ,  0.075            // 70
        , -0.444    ,  0.107            // 71
        ,  1.544    , -0.455            // 72
        ,  1.275    , -0.378            // 73
        , -1.544    , -0.455            // 74
        , -1.275    , -0.378            // 75
        ,  0.259    , -0.075            // 76
        ,  0.444    , -0.107            // 77
        , -0.259    , -0.075            // 78
        , -0.444    , -0.107            // 79
        ,  0.893    ,  0.277            // 80
        ,  1.065    ,  0.322            // 81
        , -0.893    ,  0.277            // 82
        , -1.065    ,  0.322            // 83
        ,  0.736    ,  0.228            // 84
        ,  0.594    ,   0.17            // 85
        , -0.736    ,  0.228            // 86
        , -0.594    ,   0.17            // 87
        ,  0.893    , -0.277            // 88
        ,  1.065    , -0.322            // 89
        , -0.893    , -0.277            // 90
        , -1.065    , -0.322            // 91
        ,  0.736    , -0.228            // 92
        ,  0.594    ,  -0.17            // 93
        , -0.736    , -0.228            // 94
        , -0.594    ,  -0.17            // 95
        ,  1.435    ,  0.745            // 96
        ,  1.187    ,  0.618            // 97
        , -1.435    ,  0.745            // 98
        , -1.187    ,  0.618            // 99
        ,  0.252    ,  0.194            // 100
        ,   0.37    ,   0.27            // 101
        , -0.252    ,  0.194            // 102
        ,  -0.37    ,   0.27            // 103
        ,  1.435    , -0.745            // 104
        ,  1.187    , -0.618            // 105
        , -1.435    , -0.745            // 106
        , -1.187    , -0.618            // 107
        ,  0.252    , -0.194            // 108
        ,   0.37    ,  -0.27            // 109
        , -0.252    , -0.194            // 110
        ,  -0.37    ,  -0.27            // 111
        ,  0.827    ,  0.449            // 112
        ,  0.991    ,  0.524            // 113
        , -0.827    ,  0.449            // 114
        , -0.991    ,  0.524            // 115
        ,  0.671    ,  0.386            // 116
        ,   0.52    ,  0.333            // 117
        , -0.671    ,  0.386            // 118
        ,  -0.52    ,  0.333            // 119
        ,  0.827    , -0.449            // 120
        ,  0.991    , -0.524            // 121
        , -0.827    , -0.449            // 122
        , -0.991    , -0.524            // 123
        ,  0.671    , -0.386            // 124
        ,   0.52    , -0.333            // 125
        , -0.671    , -0.386            // 126
        ,  -0.52    , -0.333            // 127
        ,  0.165    ,  1.633            // 128
        ,  0.138    ,   1.36            // 129
        , -0.165    ,  1.633            // 130
        , -0.138    ,   1.36            // 131
        ,  0.074    ,   0.09            // 132
        ,  0.074    ,  0.505            // 133
        , -0.074    ,   0.09            // 134
        , -0.074    ,  0.505            // 135
        ,  0.165    , -1.633            // 136
        ,  0.138    ,  -1.36            // 137
        , -0.165    , -1.633            // 138
        , -0.138    ,  -1.36            // 139
        ,  0.074    ,  -0.09            // 140
        ,  0.074    , -0.505            // 141
        , -0.074    ,  -0.09            // 142
        , -0.074    , -0.505            // 143
        ,  0.099    ,  0.985            // 144
        ,  0.117    ,  1.152            // 145
        , -0.099    ,  0.985            // 146
        , -0.117    ,  1.152            // 147
        ,  0.089    ,  0.829            // 148
        ,  0.089    ,  0.674            // 149
        , -0.089    ,  0.829            // 150
        , -0.089    ,  0.674            // 151
        ,  0.099    , -0.985            // 152
        ,  0.117    , -1.152            // 153
        , -0.099    , -0.985            // 154
        , -0.117    , -1.152            // 155
        ,  0.089    , -0.829            // 156
        ,  0.089    , -0.674            // 157
        , -0.089    , -0.829            // 158
        , -0.089    , -0.674            // 159
        ,  1.052    ,  1.248            // 160
        ,  0.874    ,  1.036            // 161
        , -1.052    ,  1.248            // 162
        , -0.874    ,  1.036            // 163
        ,  0.097    ,  0.245            // 164
        ,  0.196    ,  0.405            // 165
        , -0.097    ,  0.245            // 166
        , -0.196    ,  0.405            // 167
        ,  1.052    , -1.248            // 168
        ,  0.874    , -1.036            // 169
        , -1.052    , -1.248            // 170
        , -0.874    , -1.036            // 171
        ,  0.097    , -0.245            // 172
        ,  0.196    , -0.405            // 173
        , -0.097    , -0.245            // 174
        , -0.196    , -0.405            // 175
        ,  0.615    ,  0.744            // 176
        ,  0.735    ,  0.874            // 177
        , -0.615    ,  0.744            // 178
        , -0.735    ,  0.874            // 179
        ,  0.493    ,   0.63            // 180
        ,  0.362    ,  0.526            // 181
        , -0.493    ,   0.63            // 182
        , -0.362    ,  0.526            // 183
        ,  0.615    , -0.744            // 184
        ,  0.735    , -0.874            // 185
        , -0.615    , -0.744            // 186
        , -0.735    , -0.874            // 187
        ,  0.493    ,  -0.63            // 188
        ,  0.362    , -0.526            // 189
        , -0.493    ,  -0.63            // 190
        , -0.362    , -0.526            // 191
        ,  0.487    ,  1.566            // 192
        ,  0.407    ,  1.303            // 193
        , -0.487    ,  1.566            // 194
        , -0.407    ,  1.303            // 195
        ,  0.073    ,   0.09            // 196
        ,  0.088    ,    0.5            // 197
        , -0.073    ,   0.09            // 198
        , -0.088    ,    0.5            // 199
        ,  0.487    , -1.566            // 200
        ,  0.407    , -1.303            // 201
        , -0.487    , -1.566            // 202
        , -0.407    , -1.303            // 203
        ,  0.073    ,  -0.09            // 204
        ,  0.088    ,   -0.5            // 205
        , -0.073    ,  -0.09            // 206
        , -0.088    ,   -0.5            // 207
        ,  0.293    ,  0.941            // 208
        ,  0.345    ,  1.102            // 209
        , -0.293    ,  0.941            // 210
        , -0.345    ,  1.102            // 211
        ,  0.235    ,  0.795            // 212
        ,  0.167    ,  0.653            // 213
        , -0.235    ,  0.795            // 214
        , -0.167    ,  0.653            // 215
        ,  0.293    , -0.941            // 216
        ,  0.345    , -1.102            // 217
        , -0.293    , -0.941            // 218
        , -0.345    , -1.102            // 219
        ,  0.235    , -0.795            // 220
        ,  0.167    , -0.653            // 221
        , -0.235    , -0.795            // 222
        , -0.167    , -0.653            // 223
        ,  0.787    ,  1.436            // 224
        ,  0.656    ,  1.193            // 225
        , -0.787    ,  1.436            // 226
        , -0.656    ,  1.193            // 227
        ,  0.095    ,  0.245            // 228
        ,  0.187    ,  0.412            // 229
        , -0.095    ,  0.245            // 230
        , -0.187    ,  0.412            // 231
        ,  0.787    , -1.436            // 232
        ,  0.656    , -1.193            // 233
        , -0.787    , -1.436            // 234
        , -0.656    , -1.193            // 235
        ,  0.095    , -0.245            // 236
        ,  0.187    , -0.412            // 237
        , -0.095    , -0.245            // 238
        , -0.187    , -0.412            // 239
        ,  0.468    ,  0.858            // 240
        ,  0.554    ,  1.008            // 241
        , -0.468    ,  0.858            // 242
        , -0.554    ,  1.008            // 243
        ,  0.389    ,  0.714            // 244
        ,  0.311    ,  0.569            // 245
        , -0.389    ,  0.714            // 246
        , -0.311    ,  0.569            // 247
        ,  0.468    , -0.858            // 248
        ,  0.554    , -1.008            // 249
        , -0.468    , -0.858            // 250
        , -0.554    , -1.008            // 251
        ,  0.389    , -0.714            // 252
        ,  0.311    , -0.569            // 253
        , -0.389    , -0.714            // 254
        , -0.311    , -0.569            // 255
    };