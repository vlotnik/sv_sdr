    DVBS2_APSK32_8_9 : super.plane = {
            0.52    ,   0.52            // 0
        ,   0.19    ,  0.711            // 1
        ,   0.52    ,  -0.52            // 2
        ,   0.19    , -0.711            // 3
        ,  -0.52    ,   0.52            // 4
        ,  -0.19    ,  0.711            // 5
        ,  -0.52    ,  -0.52            // 6
        ,  -0.19    , -0.711            // 7
        ,  1.159    ,   0.48            // 8
        ,   0.48    ,  1.159            // 9
        ,  0.887    , -0.887            // 10
        ,      0    , -1.254            // 11
        , -0.887    ,  0.887            // 12
        ,      0    ,  1.254            // 13
        , -1.159    ,  -0.48            // 14
        ,  -0.48    , -1.159            // 15
        ,  0.711    ,   0.19            // 16
        ,  0.205    ,  0.205            // 17
        ,  0.711    ,  -0.19            // 18
        ,  0.205    , -0.205            // 19
        , -0.711    ,   0.19            // 20
        , -0.205    ,  0.205            // 21
        , -0.711    ,  -0.19            // 22
        , -0.205    , -0.205            // 23
        ,  1.254    ,      0            // 24
        ,  0.887    ,  0.887            // 25
        ,  1.159    ,  -0.48            // 26
        ,   0.48    , -1.159            // 27
        , -1.159    ,   0.48            // 28
        ,  -0.48    ,  1.159            // 29
        , -1.254    ,      0            // 30
        , -0.887    , -0.887            // 31
    };