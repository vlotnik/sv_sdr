    DVBS2_APSK16_3_4 : super.plane = {
             0.8    ,    0.8            // 0
        ,    0.8    ,   -0.8            // 1
        ,   -0.8    ,    0.8            // 2
        ,   -0.8    ,   -0.8            // 3
        ,  1.093    ,  0.293            // 4
        ,  1.093    , -0.293            // 5
        , -1.093    ,  0.293            // 6
        , -1.093    , -0.293            // 7
        ,  0.293    ,  1.093            // 8
        ,  0.293    , -1.093            // 9
        , -0.293    ,  1.093            // 10
        , -0.293    , -1.093            // 11
        ,  0.281    ,  0.281            // 12
        ,  0.281    , -0.281            // 13
        , -0.281    ,  0.281            // 14
        , -0.281    , -0.281            // 15
    };