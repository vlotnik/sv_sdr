    DVBS2_APSK16_9_10 : super.plane = {
           0.797    ,  0.797            // 0
        ,  0.797    , -0.797            // 1
        , -0.797    ,  0.797            // 2
        , -0.797    , -0.797            // 3
        ,  1.088    ,  0.292            // 4
        ,  1.088    , -0.292            // 5
        , -1.088    ,  0.292            // 6
        , -1.088    , -0.292            // 7
        ,  0.292    ,  1.088            // 8
        ,  0.292    , -1.088            // 9
        , -0.292    ,  1.088            // 10
        , -0.292    , -1.088            // 11
        ,   0.31    ,   0.31            // 12
        ,   0.31    ,  -0.31            // 13
        ,  -0.31    ,   0.31            // 14
        ,  -0.31    ,  -0.31            // 15
    };