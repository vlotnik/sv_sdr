    DVBS2X_128APSK_135_180 : super.plane = {
           0.338    ,  0.071            // 0
        ,   1.25    ,  0.427            // 1
        ,  1.317    ,  0.091            // 2
        ,  1.293    ,   0.27            // 3
        ,  0.586    ,  0.089            // 4
        ,  0.708    ,  0.187            // 5
        ,  0.948    ,  0.079            // 6
        ,  0.894    ,  0.244            // 7
        ,   0.29    ,  0.189            // 8
        ,  1.186    ,  0.582            // 9
        ,  0.996    ,  0.867            // 10
        ,  1.105    ,  0.723            // 11
        ,  0.478    ,  0.351            // 12
        ,  0.633    ,  0.368            // 13
        ,  0.726    ,  0.614            // 14
        ,  0.805    ,  0.461            // 15
        ,  0.071    ,  0.338            // 16
        ,  0.426    ,   1.25            // 17
        ,  0.092    ,  1.317            // 18
        ,   0.27    ,  1.293            // 19
        ,  0.089    ,  0.586            // 20
        ,  0.187    ,  0.708            // 21
        ,  0.079    ,  0.948            // 22
        ,  0.243    ,  0.895            // 23
        ,  0.189    ,   0.29            // 24
        ,  0.581    ,  1.186            // 25
        ,  0.866    ,  0.997            // 26
        ,  0.723    ,  1.105            // 27
        ,  0.351    ,  0.478            // 28
        ,  0.369    ,  0.633            // 29
        ,  0.614    ,  0.726            // 30
        ,  0.461    ,  0.805            // 31
        , -0.338    ,  0.071            // 32
        ,  -1.25    ,  0.427            // 33
        , -1.317    ,  0.091            // 34
        , -1.293    ,   0.27            // 35
        , -0.586    ,  0.089            // 36
        , -0.708    ,  0.187            // 37
        , -0.948    ,  0.079            // 38
        , -0.894    ,  0.244            // 39
        ,  -0.29    ,  0.189            // 40
        , -1.186    ,  0.582            // 41
        , -0.996    ,  0.867            // 42
        , -1.105    ,  0.723            // 43
        , -0.478    ,  0.351            // 44
        , -0.633    ,  0.368            // 45
        , -0.726    ,  0.614            // 46
        , -0.805    ,  0.461            // 47
        , -0.071    ,  0.338            // 48
        , -0.426    ,   1.25            // 49
        , -0.092    ,  1.317            // 50
        ,  -0.27    ,  1.293            // 51
        , -0.089    ,  0.586            // 52
        , -0.187    ,  0.708            // 53
        , -0.079    ,  0.948            // 54
        , -0.243    ,  0.895            // 55
        , -0.189    ,   0.29            // 56
        , -0.581    ,  1.186            // 57
        , -0.866    ,  0.997            // 58
        , -0.723    ,  1.105            // 59
        , -0.351    ,  0.478            // 60
        , -0.369    ,  0.633            // 61
        , -0.614    ,  0.726            // 62
        , -0.461    ,  0.805            // 63
        ,  0.338    , -0.071            // 64
        ,   1.25    , -0.427            // 65
        ,  1.317    , -0.091            // 66
        ,  1.293    ,  -0.27            // 67
        ,  0.586    , -0.089            // 68
        ,  0.708    , -0.187            // 69
        ,  0.948    , -0.079            // 70
        ,  0.894    , -0.244            // 71
        ,   0.29    , -0.189            // 72
        ,  1.186    , -0.582            // 73
        ,  0.996    , -0.867            // 74
        ,  1.105    , -0.723            // 75
        ,  0.478    , -0.351            // 76
        ,  0.633    , -0.368            // 77
        ,  0.726    , -0.614            // 78
        ,  0.805    , -0.461            // 79
        ,  0.071    , -0.338            // 80
        ,  0.426    ,  -1.25            // 81
        ,  0.092    , -1.317            // 82
        ,   0.27    , -1.293            // 83
        ,  0.089    , -0.586            // 84
        ,  0.187    , -0.708            // 85
        ,  0.079    , -0.948            // 86
        ,  0.243    , -0.895            // 87
        ,  0.189    ,  -0.29            // 88
        ,  0.581    , -1.186            // 89
        ,  0.866    , -0.997            // 90
        ,  0.723    , -1.105            // 91
        ,  0.351    , -0.478            // 92
        ,  0.369    , -0.633            // 93
        ,  0.614    , -0.726            // 94
        ,  0.461    , -0.805            // 95
        , -0.338    , -0.071            // 96
        ,  -1.25    , -0.427            // 97
        , -1.317    , -0.091            // 98
        , -1.293    ,  -0.27            // 99
        , -0.586    , -0.089            // 100
        , -0.708    , -0.187            // 101
        , -0.948    , -0.079            // 102
        , -0.894    , -0.244            // 103
        ,  -0.29    , -0.189            // 104
        , -1.186    , -0.582            // 105
        , -0.996    , -0.867            // 106
        , -1.105    , -0.723            // 107
        , -0.478    , -0.351            // 108
        , -0.633    , -0.368            // 109
        , -0.726    , -0.614            // 110
        , -0.805    , -0.461            // 111
        , -0.071    , -0.338            // 112
        , -0.426    ,  -1.25            // 113
        , -0.092    , -1.317            // 114
        ,  -0.27    , -1.293            // 115
        , -0.089    , -0.586            // 116
        , -0.187    , -0.708            // 117
        , -0.079    , -0.948            // 118
        , -0.243    , -0.895            // 119
        , -0.189    ,  -0.29            // 120
        , -0.581    , -1.186            // 121
        , -0.866    , -0.997            // 122
        , -0.723    , -1.105            // 123
        , -0.351    , -0.478            // 124
        , -0.369    , -0.633            // 125
        , -0.614    , -0.726            // 126
        , -0.461    , -0.805            // 127
    };