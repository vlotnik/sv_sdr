    QAM16_X2 : super.plane = {
           2.122    ,  2.122            // 0
        ,  2.122    ,  0.708            // 1
        ,  0.708    ,  2.122            // 2
        ,  0.708    ,  0.708            // 3
        ,  2.122    , -0.708            // 4
        ,  2.122    , -2.122            // 5
        ,  0.708    , -0.708            // 6
        ,  0.708    , -2.122            // 7
        , -0.708    ,  2.122            // 8
        , -0.708    ,  0.708            // 9
        , -2.122    ,  2.122            // 10
        , -2.122    ,  0.708            // 11
        , -0.708    , -0.708            // 12
        , -0.708    , -2.122            // 13
        , -2.122    , -0.708            // 14
        , -2.122    , -2.122            // 15
    };